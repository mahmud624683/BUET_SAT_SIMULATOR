module DFF(Q, clk, D);
input D;
input clk;
output Q;
always @(clk)
begin
  Q <= D;
end
endmodule


module c432_libar(G1gat,G4gat,G8gat,G11gat,G14gat,G17gat,G21gat,G24gat,G27gat,G30gat,G34gat,G37gat,G40gat,G43gat,G47gat,G50gat,G53gat,G56gat,G60gat,G63gat,G66gat,G69gat,G73gat,G76gat,G79gat,G82gat,G86gat,G89gat,G92gat,G95gat,G99gat,G102gat,G105gat,G108gat,G112gat,G115gat,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,G223gat,G329gat,G370gat,G421gat,G430gat,G431gat,G432gat);

input G1gat,G4gat,G8gat,G11gat,G14gat,G17gat,G21gat,G24gat,G27gat,G30gat,G34gat,G37gat,G40gat,G43gat,G47gat,G50gat,G53gat,G56gat,G60gat,G63gat,G66gat,G69gat,G73gat,G76gat,G79gat,G82gat,G86gat,G89gat,G92gat,G95gat,G99gat,G102gat,G105gat,G108gat,G112gat,G115gat,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22;
output G223gat,G329gat,G370gat,G421gat,G430gat,G431gat,G432gat;
wire G118gat,G119gat,G122gat,G123gat,G126gat,G127gat,G130gat,G131gat,G134gat,G135gat,G138gat,G139gat,G142gat,G143gat,G146gat,G147gat,G150gat,G151gat,G154gat,G157gat,CLK7,LIBAR7,RLL15,G158gat,G159gat,CLK6,LIBAR6,RLL1,G162gat,CLK5,LIBAR5,RLL20,G165gat,G168gat,G171gat,G174gat,G177gat,G180gat,G183gat,G184gat,CLK4,LIBAR4,RLL17,G185gat,G186gat,G187gat,G188gat,CLK3,LIBAR3,RLL10,G189gat,G190gat,G191gat,G192gat,G193gat,CLK2,LIBAR2,RLL11,G194gat,G195gat,G196gat,G197gat,G198gat,G1980gat,G1981gat,G199gat,G203gat,G213gat,CLK1,LIBAR1,RLL9,G224gat,RLL4,G227gat,G230gat,G233gat,G236gat,RLL14,G239gat,G242gat,RLL2,G243gat,G246gat,G247gat,G250gat,G251gat,G254gat,G255gat,G256gat,RLL16,G257gat,G258gat,G259gat,G260gat,G263gat,RLL19,G264gat,G267gat,G270gat,G273gat,G276gat,G279gat,G282gat,G285gat,RLL5,RLL18,G288gat,G289gat,RLL7,G290gat,G291gat,G292gat,G293gat,G294gat,RLL0,G295gat,G2950gat,G2951gat,G296gat,G300gat,RLL21,G301gat,G302gat,G303gat,G304gat,G305gat,G306gat,G307gat,G308gat,G309gat,G319gat,G330gat,G331gat,G332gat,G333gat,G334gat,G335gat,G336gat,G337gat,G338gat,RLL6,G339gat,G340gat,RLL13,G341gat,G342gat,G343gat,G344gat,G345gat,G346gat,RLL3,RLL22,G347gat,G348gat,G349gat,G350gat,G351gat,G352gat,G353gat,G354gat,G355gat,G356gat,G3560gat,G3561gat,G357gat,RLL12,G360gat,G371gat,G372gat,G373gat,G374gat,G375gat,G376gat,G377gat,RLL8,G378gat,G379gat,G380gat,G381gat,G386gat,G393gat,G399gat,G404gat,G407gat,G411gat,G414gat,G415gat,G4150gat,G4151gat,G416gat,G417gat,G418gat,G419gat,G420gat,G422gat,G425gat,G428gat,G429gat;

not NOT1_1 (G118gat, G1gat);
not NOT1_2 (G119gat, G4gat);
not NOT1_3 (G122gat, G11gat);
not NOT1_4 (G123gat, G17gat);
not NOT1_5 (G126gat, G24gat);
not NOT1_6 (G127gat, G30gat);
not NOT1_7 (G130gat, G37gat);
not NOT1_8 (G131gat, G43gat);
not NOT1_9 (G134gat, G50gat);
not NOT1_10 (G135gat, G56gat);
not NOT1_11 (G138gat, G63gat);
not NOT1_12 (G139gat, G69gat);
not NOT1_13 (G142gat, G76gat);
not NOT1_14 (G143gat, G82gat);
not NOT1_15 (G146gat, G89gat);
not NOT1_16 (G147gat, G95gat);
not NOT1_17 (G150gat, G102gat);
not NOT1_18 (G151gat, G108gat);
nand NAND2_19 (G154gat, G118gat, G4gat);
nor NOR2_20 (G157gat, G8gat, G119gat);
nor NOR2_21 (CLK7, G157gat, G154gat);
dff DFF2_22 (LIBAR7, CLK7, keyinput15);
xnor XNOR2_23 (RLL15, G119gat, LIBAR7);
nor NOR2_24 (G158gat, G14gat, RLL15);
nand NAND2_25 (G159gat, G122gat, G17gat);
nor NOR2_26 (CLK6, G157gat, G159gat);
dff DFF2_27 (LIBAR6, CLK6, keyinput1);
xnor XNOR2_28 (RLL1, G126gat, LIBAR6);
nand NAND2_29 (G162gat, RLL1, G30gat);
nor NOR2_30 (CLK5, G162gat, RLL1);
dff DFF2_31 (LIBAR5, CLK5, keyinput20);
xor XOR2_32 (RLL20, G130gat, LIBAR5);
nand NAND2_33 (G165gat, RLL20, G43gat);
nand NAND2_34 (G168gat, G134gat, G56gat);
nand NAND2_35 (G171gat, G138gat, G69gat);
nand NAND2_36 (G174gat, G142gat, G82gat);
nand NAND2_37 (G177gat, G146gat, G95gat);
nand NAND2_38 (G180gat, G150gat, G108gat);
nor NOR2_39 (G183gat, G21gat, G123gat);
nor NOR2_40 (G184gat, G27gat, G123gat);
nor NOR2_41 (CLK4, G162gat, G184gat);
dff DFF2_42 (LIBAR4, CLK4, keyinput17);
xnor XNOR2_43 (RLL17, G127gat, LIBAR4);
nor NOR2_44 (G185gat, G34gat, RLL17);
nor NOR2_45 (G186gat, G40gat, G127gat);
nor NOR2_46 (G187gat, G47gat, G131gat);
nor NOR2_47 (G188gat, G53gat, G131gat);
nor NOR2_48 (CLK3, G188gat, G187gat);
dff DFF2_49 (LIBAR3, CLK3, keyinput10);
xor XOR2_50 (RLL10, G135gat, LIBAR3);
nor NOR2_51 (G189gat, G60gat, RLL10);
nor NOR2_52 (G190gat, G66gat, G135gat);
nor NOR2_53 (G191gat, G73gat, G139gat);
nor NOR2_54 (G192gat, G79gat, G139gat);
nor NOR2_55 (G193gat, G86gat, G143gat);
nor NOR2_56 (CLK2, G188gat, G193gat);
dff DFF2_57 (LIBAR2, CLK2, keyinput11);
xor XOR2_58 (RLL11, G143gat, LIBAR2);
nor NOR2_59 (G194gat, G92gat, RLL11);
nor NOR2_60 (G195gat, G99gat, G147gat);
nor NOR2_61 (G196gat, G105gat, G147gat);
nor NOR2_62 (G197gat, G112gat, G151gat);
nor NOR2_63 (G198gat, G115gat, G151gat);
and AND4_64 (G1980gat, G154gat, G159gat, G162gat, G165gat);
and AND5_65 (G1981gat, G168gat, G171gat, G174gat, G177gat, G180gat);
and AND2_66 (G199gat, G1980gat, G1981gat);
not NOT1_67 (G203gat, G199gat);
not NOT1_68 (G213gat, G199gat);
nor NOR2_69 (CLK1, G213gat, G203gat);
dff DFF2_70 (LIBAR1, CLK1, keyinput9);
xor XOR2_71 (RLL9, G199gat, LIBAR1);
not NOT1_72 (G223gat, RLL9);
xor XOR2_73 (G224gat, G203gat, G154gat);
xnor XNOR2_74 (RLL4, G203gat, keyinput4);
xor XOR2_75 (G227gat, RLL4, G159gat);
xor XOR2_76 (G230gat, G203gat, G162gat);
xor XOR2_77 (G233gat, G203gat, G165gat);
xor XOR2_78 (G236gat, G203gat, G168gat);
xnor XNOR2_79 (RLL14, G203gat, keyinput14);
xor XOR2_80 (G239gat, RLL14, G171gat);
nand NAND2_81 (G242gat, G1gat, G213gat);
xor XOR2_82 (RLL2, G203gat, keyinput2);
xor XOR2_83 (G243gat, RLL2, G174gat);
nand NAND2_84 (G246gat, G213gat, G11gat);
xor XOR2_85 (G247gat, G203gat, G177gat);
nand NAND2_86 (G250gat, G213gat, G24gat);
xor XOR2_87 (G251gat, G203gat, G180gat);
nand NAND2_88 (G254gat, G213gat, G37gat);
nand NAND2_89 (G255gat, G213gat, G50gat);
nand NAND2_90 (G256gat, G213gat, G63gat);
xor XOR2_91 (RLL16, G213gat, keyinput16);
nand NAND2_92 (G257gat, RLL16, G76gat);
nand NAND2_93 (G258gat, G213gat, G89gat);
nand NAND2_94 (G259gat, G213gat, G102gat);
nand NAND2_95 (G260gat, G224gat, G157gat);
nand NAND2_96 (G263gat, G224gat, G158gat);
xnor XNOR2_97 (RLL19, G227gat, keyinput19);
nand NAND2_98 (G264gat, RLL19, G183gat);
nand NAND2_99 (G267gat, G230gat, G185gat);
nand NAND2_100 (G270gat, G233gat, G187gat);
nand NAND2_101 (G273gat, G236gat, G189gat);
nand NAND2_102 (G276gat, G239gat, G191gat);
nand NAND2_103 (G279gat, G243gat, G193gat);
nand NAND2_104 (G282gat, G247gat, G195gat);
nand NAND2_105 (G285gat, G251gat, G197gat);
xor XOR2_106 (RLL5, G227gat, keyinput5);
xor XOR2_107 (RLL18, RLL5, keyinput18);
nand NAND2_108 (G288gat, RLL18, G184gat);
nand NAND2_109 (G289gat, G230gat, G186gat);
xor XOR2_110 (RLL7, G233gat, keyinput7);
nand NAND2_111 (G290gat, RLL7, G188gat);
nand NAND2_112 (G291gat, G236gat, G190gat);
nand NAND2_113 (G292gat, G239gat, G192gat);
nand NAND2_114 (G293gat, G243gat, G194gat);
nand NAND2_115 (G294gat, G247gat, G196gat);
xor XOR2_116 (RLL0, G251gat, keyinput0);
nand NAND2_117 (G295gat, RLL0, G198gat);
and AND4_118 (G2950gat, G260gat, G264gat, G267gat, G270gat);
and AND5_119 (G2951gat, G273gat, G276gat, G279gat, G282gat, G285gat);
and AND2_120 (G296gat, G2950gat, G2951gat);
not NOT1_121 (G300gat, G263gat);
xnor XNOR2_122 (RLL21, G288gat, keyinput21);
not NOT1_123 (G301gat, RLL21);
not NOT1_124 (G302gat, G289gat);
not NOT1_125 (G303gat, G290gat);
not NOT1_126 (G304gat, G291gat);
not NOT1_127 (G305gat, G292gat);
not NOT1_128 (G306gat, G293gat);
not NOT1_129 (G307gat, G294gat);
not NOT1_130 (G308gat, G295gat);
not NOT1_131 (G309gat, G296gat);
not NOT1_132 (G319gat, G296gat);
not NOT1_133 (G329gat, G296gat);
xor XOR2_134 (G330gat, G309gat, G260gat);
xor XOR2_135 (G331gat, G309gat, G264gat);
xor XOR2_136 (G332gat, G309gat, G267gat);
xor XOR2_137 (G333gat, G309gat, G270gat);
nand NAND2_138 (G334gat, G8gat, G319gat);
xor XOR2_139 (G335gat, G309gat, G273gat);
nand NAND2_140 (G336gat, G319gat, G21gat);
xor XOR2_141 (G337gat, G309gat, G276gat);
nand NAND2_142 (G338gat, G319gat, G34gat);
xnor XNOR2_143 (RLL6, G309gat, keyinput6);
xor XOR2_144 (G339gat, RLL6, G279gat);
nand NAND2_145 (G340gat, G319gat, G47gat);
xnor XNOR2_146 (RLL13, G309gat, keyinput13);
xor XOR2_147 (G341gat, RLL13, G282gat);
nand NAND2_148 (G342gat, G319gat, G60gat);
xor XOR2_149 (G343gat, G309gat, G285gat);
nand NAND2_150 (G344gat, G319gat, G73gat);
nand NAND2_151 (G345gat, G319gat, G86gat);
nand NAND2_152 (G346gat, G319gat, G99gat);
xnor XNOR2_153 (RLL3, G319gat, keyinput3);
xnor XNOR2_154 (RLL22, RLL3, keyinput22);
nand NAND2_155 (G347gat, RLL22, G112gat);
nand NAND2_156 (G348gat, G330gat, G300gat);
nand NAND2_157 (G349gat, G331gat, G301gat);
nand NAND2_158 (G350gat, G332gat, G302gat);
nand NAND2_159 (G351gat, G333gat, G303gat);
nand NAND2_160 (G352gat, G335gat, G304gat);
nand NAND2_161 (G353gat, G337gat, G305gat);
nand NAND2_162 (G354gat, G339gat, G306gat);
nand NAND2_163 (G355gat, G341gat, G307gat);
nand NAND2_164 (G356gat, G343gat, G308gat);
and AND4_165 (G3560gat, G348gat, G349gat, G350gat, G351gat);
and AND5_166 (G3561gat, G352gat, G353gat, G354gat, G355gat, G356gat);
and AND2_167 (G357gat, G3560gat, G3561gat);
xnor XNOR2_168 (RLL12, G357gat, keyinput12);
not NOT1_169 (G360gat, RLL12);
not NOT1_170 (G370gat, G357gat);
nand NAND2_171 (G371gat, G14gat, G360gat);
nand NAND2_172 (G372gat, G360gat, G27gat);
nand NAND2_173 (G373gat, G360gat, G40gat);
nand NAND2_174 (G374gat, G360gat, G53gat);
nand NAND2_175 (G375gat, G360gat, G66gat);
nand NAND2_176 (G376gat, G360gat, G79gat);
nand NAND2_177 (G377gat, G360gat, G92gat);
xor XOR2_178 (RLL8, G360gat, keyinput8);
nand NAND2_179 (G378gat, RLL8, G105gat);
nand NAND2_180 (G379gat, G360gat, G115gat);
nand NAND4_181 (G380gat, G4gat, G242gat, G334gat, G371gat);
nand NAND4_182 (G381gat, G246gat, G336gat, G372gat, G17gat);
nand NAND4_183 (G386gat, G250gat, G338gat, G373gat, G30gat);
nand NAND4_184 (G393gat, G254gat, G340gat, G374gat, G43gat);
nand NAND4_185 (G399gat, G255gat, G342gat, G375gat, G56gat);
nand NAND4_186 (G404gat, G256gat, G344gat, G376gat, G69gat);
nand NAND4_187 (G407gat, G257gat, G345gat, G377gat, G82gat);
nand NAND4_188 (G411gat, G258gat, G346gat, G378gat, G95gat);
nand NAND4_189 (G414gat, G259gat, G347gat, G379gat, G108gat);
not NOT1_190 (G415gat, G380gat);
and AND4_191 (G4150gat, G381gat, G386gat, G393gat, G399gat);
and AND4_192 (G4151gat, G404gat, G407gat, G411gat, G414gat);
and AND2_193 (G416gat, G4150gat, G4151gat);
not NOT1_194 (G417gat, G393gat);
not NOT1_195 (G418gat, G404gat);
not NOT1_196 (G419gat, G407gat);
not NOT1_197 (G420gat, G411gat);
nor NOR2_198 (G421gat, G415gat, G416gat);
nand NAND2_199 (G422gat, G386gat, G417gat);
nand NAND4_200 (G425gat, G386gat, G393gat, G418gat, G399gat);
nand NAND3_201 (G428gat, G399gat, G393gat, G419gat);
nand NAND4_202 (G429gat, G386gat, G393gat, G407gat, G420gat);
nand NAND4_203 (G430gat, G381gat, G386gat, G422gat, G399gat);
nand NAND4_204 (G431gat, G381gat, G386gat, G425gat, G428gat);
nand NAND4_205 (G432gat, G381gat, G422gat, G425gat, G429gat);

endmodule