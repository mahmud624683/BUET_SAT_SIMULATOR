module c1908_rll_8k(G1gat,G4gat,G7gat,G10gat,G13gat,G16gat,G19gat,G22gat,G25gat,G28gat,G31gat,G34gat,G37gat,G40gat,G43gat,G46gat,G49gat,G53gat,G56gat,G60gat,G63gat,G66gat,G69gat,G72gat,G76gat,G79gat,G82gat,G85gat,G88gat,G91gat,G94gat,G99gat,G104gat,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,G2753gat,G2754gat,G2755gat,G2756gat,G2762gat,G2767gat,G2768gat,G2779gat,G2780gat,G2781gat,G2782gat,G2783gat,G2784gat,G2785gat,G2786gat,G2787gat,G2811gat,G2886gat,G2887gat,G2888gat,G2889gat,G2890gat,G2891gat,G2892gat,G2899gat);

input G1gat,G4gat,G7gat,G10gat,G13gat,G16gat,G19gat,G22gat,G25gat,G28gat,G31gat,G34gat,G37gat,G40gat,G43gat,G46gat,G49gat,G53gat,G56gat,G60gat,G63gat,G66gat,G69gat,G72gat,G76gat,G79gat,G82gat,G85gat,G88gat,G91gat,G94gat,G99gat,G104gat,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7;
output G2753gat,G2754gat,G2755gat,G2756gat,G2762gat,G2767gat,G2768gat,G2779gat,G2780gat,G2781gat,G2782gat,G2783gat,G2784gat,G2785gat,G2786gat,G2787gat,G2811gat,G2886gat,G2887gat,G2888gat,G2889gat,G2890gat,G2891gat,G2892gat,G2899gat;
wire G190gat_enc,G190gat,G194gat_enc,G194gat,G197gat_enc,G197gat,G201gat,G206gat_enc,G206gat,G209gat_enc,G209gat,G212gat_enc,G212gat,G216gat_enc,G216gat,G220gat_enc,G220gat,G225gat,G229gat,G232gat,G235gat,G239gat,G243gat,G247gat,G251gat,G252gat,G253gat,G256gat,G263gat,G266gat,G269gat,G272gat,G275gat,G276gat,G277gat,G280gat,G290gat,G300gat,G306gat,G313gat,G319gat,G338gat,G534gat,G535gat,G536gat,G537gat,G538gat,G539gat,G540gat,G541gat,G542gat,G543gat,G544gat,G545gat,G546gat,G547gat,G548gat,G549gat,G550gat,G551gat,G552gat,G553gat,G554gat,G555gat,G574gat,G586gat,G592gat,G601gat,G602gat,G603gat,G608gat,G612gat,G643gat,G655gat,G682gat,G685gat,G724gat,G886gat,G887gat,G888gat,G889gat,G890gat,G891gat,G892gat,G893gat,G894gat,G895gat,G896gat,G897gat,G898gat,G899gat,G903gat,G907gat,G910gat,G913gat,G914gat,G915gat,G916gat,G917gat,G918gat,G919gat,G920gat,G921gat,G922gat,G923gat,G926gat,G938gat,G942gat,G946gat,G950gat,G954gat,G958gat,G968gat,G972gat,G976gat,G980gat,G984gat,G988gat,G989gat,G990gat,G991gat,G992gat,G993gat,G997gat,G1001gat,G1002gat,G1003gat,G1004gat,G1005gat,G1006gat,G1007gat,G1008gat,G1009gat,G1054gat,G1055gat,G1063gat,G1064gat,G1067gat,G1068gat,G1119gat,G1120gat,G1121gat,G1122gat,G1128gat,G1129gat,G1130gat,G1131gat,G1132gat,G1133gat,G1148gat,G1149gat,G1150gat,G1151gat,G1152gat,G1153gat,G1154gat,G1155gat,G1156gat,G1157gat,G1158gat,G1159gat,G1160gat,G1161gat,G1162gat,G1163gat,G1167gat,G1171gat,G1188gat,G1205gat,G1206gat,G1207gat,G1208gat,G1209gat,G1210gat,G1211gat,G1212gat,G1213gat,G1214gat,G1215gat,G1216gat,G1217gat,G1218gat,G1219gat,G1220gat,G1221gat,G1222gat,G1223gat,G1224gat,G1225gat,G1226gat,G1227gat,G1228gat,G1229gat,G1230gat,G1231gat,G1232gat,G1235gat,G1238gat,G1239gat,G1240gat,G1241gat,G1242gat,G1243gat,G1246gat,G1249gat,G1264gat,G1267gat,G1309gat,G1310gat,G1311gat,G1312gat,G1313gat,G1314gat,G1315gat,G1316gat,G1317gat,G1318gat,G1319gat,G1322gat,G1327gat,G1328gat,G1334gat,G1344gat,G1345gat,G1346gat,G1348gat,G1349gat,G1350gat,G1351gat,G1352gat,G1355gat,G1358gat,G1361gat,G1364gat,G1367gat,G1370gat,G1373gat,G1376gat,G1379gat,G1383gat,G1386gat,G1387gat,G1388gat,G1389gat,G1390gat,G1393gat,G1396gat,G1397gat,G1398gat,G1399gat,G1409gat,G1412gat,G1413gat,G1433gat,G1434gat,G1438gat,G1439gat,G1440gat,G1443gat,G1444gat,G1445gat,G1446gat,G1447gat,G1448gat,G1451gat,G1452gat,G1453gat,G1454gat,G1455gat,G1456gat,G1457gat,G1458gat,G1459gat,G1460gat,G1461gat,G1462gat,G1463gat,G1464gat,G1468gat,G1469gat,G1470gat,G1471gat,G1472gat,G1475gat,G1476gat,G1478gat,G1481gat,G1484gat,G1487gat,G1488gat,G1489gat,G1490gat,G1491gat,G1492gat,G1493gat,G1494gat,G1495gat,G1496gat,G1498gat,G1499gat,G1500gat,G1501gat,G1504gat,G1510gat,G1513gat,G1514gat,G1517gat,G1520gat,G1521gat,G1522gat,G1526gat,G1527gat,G1528gat,G1529gat,G1530gat,G1531gat,G1532gat,G1534gat,G1537gat,G1540gat,G1546gat,G1554gat,G1557gat,G1561gat,G1567gat,G1568gat,G1569gat,G1571gat,G1576gat,G1591gat,G1593gat,G1594gat,G1595gat,G1596gat,G1635gat,G1636gat,G1638gat,G1639gat,G1671gat,G1672gat,G1675gat,G1677gat,G1678gat,G1679gat,G1680gat,G1681gat,G1682gat,G1683gat,G1685gat,G1688gat,G1706gat,G1707gat,G1708gat,G1709gat,G1710gat,G1711gat,G1712gat,G1713gat,G1720gat,G1721gat,G1723gat,G1727gat,G1728gat,G1730gat,G1740gat,G1741gat,G1742gat,G1746gat,G1747gat,G1748gat,G1751gat,G1759gat,G1761gat,G1762gat,G1763gat,G1764gat,G1768gat,G1769gat,G1772gat,G1773gat,G1774gat,G1777gat,G1783gat,G1784gat,G1785gat,G1786gat,G1787gat,G1788gat,G1791gat,G1792gat,G1795gat,G1796gat,G1798gat,G1801gat,G1802gat,G1807gat,G1808gat,G1809gat,G1810gat,G1812gat,G1815gat,G1821gat,G1822gat,G1823gat,G1824gat,G1825gat,G1826gat,G1827gat,G1830gat,G1837gat,G1838gat,G1841gat,G1848gat,G1849gat,G1850gat,G1852gat,G1855gat,G1856gat,G1857gat,G1858gat,G1864gat,G1865gat,G1875gat,G1878gat,G1879gat,G1882gat,G1883gat,G1884gat,G1885gat,G1889gat,G1895gat,G1896gat,G1897gat,G1898gat,G1910gat,G1911gat,G1912gat,G1913gat,G1915gat,G1919gat,G1920gat,G1921gat,G1922gat,G1923gat,G1924gat,G1933gat,G1936gat,G1937gat,G1938gat,G1941gat,G1942gat,G1947gat,G1961gat,G1965gat,G1968gat,G1975gat,G1976gat,G1977gat,G1978gat,G1979gat,G1980gat,G1985gat,G1987gat,G1999gat,G2000gat,G2002gat,G2003gat,G2004gat,G2005gat,G2006gat,G2007gat,G2008gat,G2009gat,G2012gat,G2013gat,G2014gat,G2015gat,G2016gat,G2018gat,G2019gat,G2020gat,G2021gat,G2022gat,G2023gat,G2024gat,G2025gat,G2026gat,G2027gat,G2030gat,G2036gat,G2037gat,G2038gat,G2039gat,G2040gat,G2041gat,G2042gat,G2047gat,G2052gat,G2055gat,G2060gat,G2061gat,G2062gat,G2067gat,G2068gat,G2076gat,G2077gat,G2078gat,G2081gat,G2086gat,G2104gat,G2119gat,G2129gat,G2143gat,G2214gat,G2215gat,G2216gat,G2217gat,G2222gat,G2223gat,G2224gat,G2225gat,G2226gat,G2227gat,G2228gat,G2229gat,G2230gat,G2231gat,G2232gat,G2233gat,G2234gat,G2235gat,G2236gat,G2237gat,G2240gat,G2241gat,G2244gat,G2245gat,G2250gat,G2253gat,G2256gat,G2257gat,G2263gat,G2266gat,G2269gat,G2272gat,G2273gat,G2274gat,G2279gat,G2340gat,G2353gat,G2361gat,G2375gat,G2384gat,G2385gat,G2386gat,G2426gat,G2427gat,G2537gat,G2540gat,G2543gat,G2546gat,G2549gat,G2552gat,G2555gat,G2558gat,G2561gat,G2564gat,G2567gat,G2570gat,G2573gat,G2576gat,G2594gat,G2597gat,G2600gat,G2603gat,G2606gat,G2611gat,G2614gat,G2617gat,G2620gat,G2627gat,G2628gat,G2629gat,G2630gat,G2631gat,G2632gat,G2633gat,G2634gat,G2639gat,G2642gat,G2645gat,G2648gat,G2651gat,G2655gat,G2658gat,G2661gat,G2664gat,G2669gat,G2670gat,G2671gat,G2672gat,G2673gat,G2674gat,G2675gat,G2676gat,G2682gat,G2683gat,G2688gat,G2689gat,G2690gat,G2691gat,G2692gat,G2693gat,G2710gat,G2720gat,G2721gat,G2722gat,G2723gat,G2724gat,G2725gat,G2726gat,G2727gat,G2728gat,G2729gat,G2730gat,G2731gat,G2732gat,G2733gat,G2734gat,G2735gat,G2736gat,G2737gat,G2738gat,G2739gat,G2740gat,G2741gat,G2742gat,G2743gat,G2744gat,G27440gat,G27441gat,G2745gat,G27450gat,G27451gat,G2746gat,G27460gat,G27461gat,G2747gat,G27470gat,G27471gat,G2750gat,G2757gat,G2758gat,G2759gat,G2760gat,G2761gat,G2763gat,G2764gat,G2765gat,G2766gat,G2773gat,G2776gat,G2788gat,G2789gat,G2800gat,G2807gat,G2808gat,G2809gat,G2810gat,G2812gat,G2815gat,G2818gat,G2821gat,G2824gat,G2827gat,G2828gat,G2829gat,G2843gat,G2846gat,G2850gat,G2851gat,G2852gat,G2853gat,G2854gat,G2857gat,G2858gat,G2859gat,G2860gat,G2861gat,G2862gat,G2863gat,G2866gat,G2867gat,G2868gat,G2869gat,G2870gat,G2871gat,G2872gat,G2873gat,G2874gat,G2875gat,G2876gat,G2877gat,G2878gat,G2879gat,G2880gat,G2881gat,G2882gat,G2883gat,G2895gat,G2896gat,G2897gat,G2898gat;

not NOT1_1 (G190gat_enc, G1gat);
xnor XNOR2_2 (G190gat, keyinput0, G190gat_enc);
not NOT1_3 (G194gat_enc, G4gat);
xor XOR2_4 (G194gat, keyinput1, G194gat_enc);
not NOT1_5 (G197gat_enc, G7gat);
xnor XNOR2_6 (G197gat, keyinput2, G197gat_enc);
not NOT1_7 (G201gat, G10gat);
not NOT1_8 (G206gat_enc, G13gat);
xnor XNOR2_9 (G206gat, keyinput3, G206gat_enc);
not NOT1_10 (G209gat_enc, G16gat);
xor XOR2_11 (G209gat, keyinput4, G209gat_enc);
not NOT1_12 (G212gat_enc, G19gat);
xor XOR2_13 (G212gat, keyinput5, G212gat_enc);
not NOT1_14 (G216gat_enc, G22gat);
xnor XNOR2_15 (G216gat, keyinput6, G216gat_enc);
not NOT1_16 (G220gat_enc, G25gat);
xor XOR2_17 (G220gat, keyinput7, G220gat_enc);
not NOT1_18 (G225gat, G28gat);
not NOT1_19 (G229gat, G31gat);
not NOT1_20 (G232gat, G34gat);
not NOT1_21 (G235gat, G37gat);
not NOT1_22 (G239gat, G40gat);
not NOT1_23 (G243gat, G43gat);
not NOT1_24 (G247gat, G46gat);
nand NAND2_25 (G251gat, G63gat, G88gat);
nand NAND2_26 (G252gat, G66gat, G91gat);
not NOT1_27 (G253gat, G72gat);
not NOT1_28 (G256gat, G72gat);
not NOT1_29 (G263gat, G76gat);
not NOT1_30 (G266gat, G79gat);
not NOT1_31 (G269gat, G82gat);
not NOT1_32 (G272gat, G85gat);
not NOT1_33 (G275gat, G104gat);
not NOT1_34 (G276gat, G104gat);
not NOT1_35 (G277gat, G88gat);
not NOT1_36 (G280gat, G91gat);
not NOT1_37 (G290gat, G94gat);
not NOT1_38 (G300gat, G94gat);
not NOT1_39 (G306gat, G99gat);
not NOT1_40 (G313gat, G99gat);
not NOT1_41 (G319gat, G104gat);
not NOT1_42 (G338gat, G104gat);
not NOT1_43 (G534gat, G343gat);
not NOT1_44 (G535gat, G346gat);
not NOT1_45 (G536gat, G349gat);
not NOT1_46 (G537gat, G352gat);
not NOT1_47 (G538gat, G355gat);
not NOT1_48 (G539gat, G358gat);
not NOT1_49 (G540gat, G361gat);
not NOT1_50 (G541gat, G364gat);
not NOT1_51 (G542gat, G367gat);
not NOT1_52 (G543gat, G370gat);
not NOT1_53 (G544gat, G373gat);
not NOT1_54 (G545gat, G376gat);
not NOT1_55 (G546gat, G379gat);
not NOT1_56 (G547gat, G382gat);
not NOT1_57 (G548gat, G385gat);
not NOT1_58 (G549gat, G388gat);
nand NAND2_59 (G550gat, G306gat, G331gat);
nand NAND2_60 (G551gat, G306gat, G331gat);
nand NAND2_61 (G552gat, G306gat, G331gat);
nand NAND2_62 (G553gat, G306gat, G331gat);
nand NAND2_63 (G554gat, G306gat, G331gat);
nand NAND2_64 (G555gat, G306gat, G331gat);
and AND2_65 (G574gat, G63gat, G319gat);
and AND2_66 (G586gat, G66gat, G319gat);
and AND3_67 (G592gat, G49gat, G253gat, G319gat);
nand NAND2_68 (G601gat, G326gat, G277gat);
nand NAND2_69 (G602gat, G326gat, G280gat);
nand NAND2_70 (G603gat, G260gat, G72gat);
nand NAND2_71 (G608gat, G260gat, G300gat);
nand NAND2_72 (G612gat, G256gat, G300gat);
and AND3_73 (G643gat, G56gat, G257gat, G319gat);
and AND3_74 (G655gat, G60gat, G257gat, G319gat);
and AND2_75 (G682gat, G251gat, G316gat);
and AND2_76 (G685gat, G252gat, G316gat);
and AND3_77 (G724gat, G53gat, G253gat, G319gat);
not NOT1_78 (G886gat, G682gat);
not NOT1_79 (G887gat, G685gat);
not NOT1_80 (G888gat, G616gat);
not NOT1_81 (G889gat, G619gat);
not NOT1_82 (G890gat, G622gat);
not NOT1_83 (G891gat, G625gat);
not NOT1_84 (G892gat, G631gat);
not NOT1_85 (G893gat, G643gat);
not NOT1_86 (G894gat, G649gat);
not NOT1_87 (G895gat, G652gat);
not NOT1_88 (G896gat, G655gat);
and AND2_89 (G897gat, G49gat, G612gat);
and AND2_90 (G898gat, G56gat, G608gat);
nand NAND2_91 (G899gat, G53gat, G612gat);
nand NAND2_92 (G903gat, G60gat, G608gat);
nand NAND2_93 (G907gat, G49gat, G612gat);
nand NAND2_94 (G910gat, G56gat, G608gat);
not NOT1_95 (G913gat, G661gat);
not NOT1_96 (G914gat, G658gat);
not NOT1_97 (G915gat, G667gat);
not NOT1_98 (G916gat, G664gat);
not NOT1_99 (G917gat, G673gat);
not NOT1_100 (G918gat, G670gat);
not NOT1_101 (G919gat, G679gat);
not NOT1_102 (G920gat, G676gat);
nand NAND4_103 (G921gat, G277gat, G297gat, G326gat, G603gat);
nand NAND4_104 (G922gat, G280gat, G297gat, G326gat, G603gat);
nand NAND3_105 (G923gat, G303gat, G338gat, G603gat);
and AND3_106 (G926gat, G303gat, G338gat, G603gat);
not NOT1_107 (G938gat, G688gat);
not NOT1_108 (G942gat, G691gat);
not NOT1_109 (G946gat, G694gat);
not NOT1_110 (G950gat, G697gat);
not NOT1_111 (G954gat, G700gat);
not NOT1_112 (G958gat, G703gat);
not NOT1_113 (G968gat, G706gat);
not NOT1_114 (G972gat, G709gat);
not NOT1_115 (G976gat, G712gat);
not NOT1_116 (G980gat, G715gat);
not NOT1_117 (G984gat, G628gat);
not NOT1_118 (G988gat, G718gat);
not NOT1_119 (G989gat, G721gat);
not NOT1_120 (G990gat, G634gat);
not NOT1_121 (G991gat, G724gat);
not NOT1_122 (G992gat, G727gat);
not NOT1_123 (G993gat, G637gat);
not NOT1_124 (G997gat, G730gat);
not NOT1_125 (G1001gat, G733gat);
not NOT1_126 (G1002gat, G736gat);
not NOT1_127 (G1003gat, G739gat);
not NOT1_128 (G1004gat, G640gat);
not NOT1_129 (G1005gat, G742gat);
not NOT1_130 (G1006gat, G745gat);
not NOT1_131 (G1007gat, G646gat);
not NOT1_132 (G1008gat, G748gat);
not NOT1_133 (G1009gat, G751gat);
nand NAND2_134 (G1054gat, G619gat, G888gat);
nand NAND2_135 (G1055gat, G616gat, G889gat);
nand NAND2_136 (G1063gat, G625gat, G890gat);
nand NAND2_137 (G1064gat, G622gat, G891gat);
nand NAND2_138 (G1067gat, G655gat, G895gat);
nand NAND2_139 (G1068gat, G652gat, G896gat);
nand NAND2_140 (G1119gat, G721gat, G988gat);
nand NAND2_141 (G1120gat, G718gat, G989gat);
nand NAND2_142 (G1121gat, G727gat, G991gat);
nand NAND2_143 (G1122gat, G724gat, G992gat);
nand NAND2_144 (G1128gat, G739gat, G1002gat);
nand NAND2_145 (G1129gat, G736gat, G1003gat);
nand NAND2_146 (G1130gat, G745gat, G1005gat);
nand NAND2_147 (G1131gat, G742gat, G1006gat);
nand NAND2_148 (G1132gat, G751gat, G1008gat);
nand NAND2_149 (G1133gat, G748gat, G1009gat);
not NOT1_150 (G1148gat, G939gat);
not NOT1_151 (G1149gat, G935gat);
nand NAND2_152 (G1150gat, G1054gat, G1055gat);
not NOT1_153 (G1151gat, G943gat);
not NOT1_154 (G1152gat, G947gat);
not NOT1_155 (G1153gat, G955gat);
not NOT1_156 (G1154gat, G951gat);
not NOT1_157 (G1155gat, G962gat);
not NOT1_158 (G1156gat, G969gat);
not NOT1_159 (G1157gat, G977gat);
nand NAND2_160 (G1158gat, G1063gat, G1064gat);
not NOT1_161 (G1159gat, G985gat);
nand NAND2_162 (G1160gat, G985gat, G892gat);
not NOT1_163 (G1161gat, G998gat);
nand NAND2_164 (G1162gat, G1067gat, G1068gat);
not NOT1_165 (G1163gat, G899gat);
not NOT1_166 (G1167gat, G903gat);
nand NAND2_167 (G1171gat, G921gat, G923gat);
nand NAND2_168 (G1188gat, G922gat, G923gat);
not NOT1_169 (G1205gat, G1010gat);
nand NAND2_170 (G1206gat, G1010gat, G938gat);
not NOT1_171 (G1207gat, G1013gat);
nand NAND2_172 (G1208gat, G1013gat, G942gat);
not NOT1_173 (G1209gat, G1016gat);
nand NAND2_174 (G1210gat, G1016gat, G946gat);
not NOT1_175 (G1211gat, G1019gat);
nand NAND2_176 (G1212gat, G1019gat, G950gat);
not NOT1_177 (G1213gat, G1022gat);
nand NAND2_178 (G1214gat, G1022gat, G954gat);
not NOT1_179 (G1215gat, G1025gat);
nand NAND2_180 (G1216gat, G1025gat, G958gat);
not NOT1_181 (G1217gat, G1028gat);
not NOT1_182 (G1218gat, G959gat);
not NOT1_183 (G1219gat, G1031gat);
not NOT1_184 (G1220gat, G1034gat);
nand NAND2_185 (G1221gat, G1034gat, G968gat);
not NOT1_186 (G1222gat, G965gat);
not NOT1_187 (G1223gat, G1037gat);
nand NAND2_188 (G1224gat, G1037gat, G972gat);
not NOT1_189 (G1225gat, G1040gat);
nand NAND2_190 (G1226gat, G1040gat, G976gat);
not NOT1_191 (G1227gat, G973gat);
not NOT1_192 (G1228gat, G1043gat);
nand NAND2_193 (G1229gat, G1043gat, G980gat);
not NOT1_194 (G1230gat, G981gat);
nand NAND2_195 (G1231gat, G981gat, G984gat);
nand NAND2_196 (G1232gat, G1119gat, G1120gat);
nand NAND2_197 (G1235gat, G1121gat, G1122gat);
not NOT1_198 (G1238gat, G1046gat);
nand NAND2_199 (G1239gat, G1046gat, G997gat);
not NOT1_200 (G1240gat, G994gat);
not NOT1_201 (G1241gat, G1049gat);
nand NAND2_202 (G1242gat, G1049gat, G1001gat);
nand NAND2_203 (G1243gat, G1128gat, G1129gat);
nand NAND2_204 (G1246gat, G1130gat, G1131gat);
nand NAND2_205 (G1249gat, G1132gat, G1133gat);
not NOT1_206 (G1264gat, G1150gat);
nand NAND2_207 (G1267gat, G631gat, G1159gat);
nand NAND2_208 (G1309gat, G688gat, G1205gat);
nand NAND2_209 (G1310gat, G691gat, G1207gat);
nand NAND2_210 (G1311gat, G694gat, G1209gat);
nand NAND2_211 (G1312gat, G697gat, G1211gat);
nand NAND2_212 (G1313gat, G700gat, G1213gat);
nand NAND2_213 (G1314gat, G703gat, G1215gat);
nand NAND2_214 (G1315gat, G706gat, G1220gat);
nand NAND2_215 (G1316gat, G709gat, G1223gat);
nand NAND2_216 (G1317gat, G712gat, G1225gat);
nand NAND2_217 (G1318gat, G715gat, G1228gat);
not NOT1_218 (G1319gat, G1158gat);
nand NAND2_219 (G1322gat, G628gat, G1230gat);
nand NAND2_220 (G1327gat, G730gat, G1238gat);
nand NAND2_221 (G1328gat, G733gat, G1241gat);
not NOT1_222 (G1334gat, G1162gat);
nand NAND2_223 (G1344gat, G1267gat, G1160gat);
nand NAND2_224 (G1345gat, G1249gat, G894gat);
not NOT1_225 (G1346gat, G1249gat);
not NOT1_226 (G1348gat, G1255gat);
not NOT1_227 (G1349gat, G1252gat);
not NOT1_228 (G1350gat, G1261gat);
not NOT1_229 (G1351gat, G1258gat);
nand NAND2_230 (G1352gat, G1309gat, G1206gat);
nand NAND2_231 (G1355gat, G1310gat, G1208gat);
nand NAND2_232 (G1358gat, G1311gat, G1210gat);
nand NAND2_233 (G1361gat, G1312gat, G1212gat);
nand NAND2_234 (G1364gat, G1313gat, G1214gat);
nand NAND2_235 (G1367gat, G1314gat, G1216gat);
nand NAND2_236 (G1370gat, G1315gat, G1221gat);
nand NAND2_237 (G1373gat, G1316gat, G1224gat);
nand NAND2_238 (G1376gat, G1317gat, G1226gat);
nand NAND2_239 (G1379gat, G1318gat, G1229gat);
nand NAND2_240 (G1383gat, G1322gat, G1231gat);
not NOT1_241 (G1386gat, G1232gat);
nand NAND2_242 (G1387gat, G1232gat, G990gat);
not NOT1_243 (G1388gat, G1235gat);
nand NAND2_244 (G1389gat, G1235gat, G993gat);
nand NAND2_245 (G1390gat, G1327gat, G1239gat);
nand NAND2_246 (G1393gat, G1328gat, G1242gat);
not NOT1_247 (G1396gat, G1243gat);
nand NAND2_248 (G1397gat, G1243gat, G1004gat);
not NOT1_249 (G1398gat, G1246gat);
nand NAND2_250 (G1399gat, G1246gat, G1007gat);
not NOT1_251 (G1409gat, G1319gat);
nand NAND2_252 (G1412gat, G649gat, G1346gat);
not NOT1_253 (G1413gat, G1334gat);
nand NAND2_254 (G1433gat, G634gat, G1386gat);
nand NAND2_255 (G1434gat, G637gat, G1388gat);
nand NAND2_256 (G1438gat, G640gat, G1396gat);
nand NAND2_257 (G1439gat, G646gat, G1398gat);
not NOT1_258 (G1440gat, G1344gat);
nand NAND2_259 (G1443gat, G1355gat, G1148gat);
not NOT1_260 (G1444gat, G1355gat);
nand NAND2_261 (G1445gat, G1352gat, G1149gat);
not NOT1_262 (G1446gat, G1352gat);
nand NAND2_263 (G1447gat, G1358gat, G1151gat);
not NOT1_264 (G1448gat, G1358gat);
nand NAND2_265 (G1451gat, G1361gat, G1152gat);
not NOT1_266 (G1452gat, G1361gat);
nand NAND2_267 (G1453gat, G1367gat, G1153gat);
not NOT1_268 (G1454gat, G1367gat);
nand NAND2_269 (G1455gat, G1364gat, G1154gat);
not NOT1_270 (G1456gat, G1364gat);
nand NAND2_271 (G1457gat, G1373gat, G1156gat);
not NOT1_272 (G1458gat, G1373gat);
nand NAND2_273 (G1459gat, G1379gat, G1157gat);
not NOT1_274 (G1460gat, G1379gat);
not NOT1_275 (G1461gat, G1383gat);
nand NAND2_276 (G1462gat, G1393gat, G1161gat);
not NOT1_277 (G1463gat, G1393gat);
nand NAND2_278 (G1464gat, G1345gat, G1412gat);
not NOT1_279 (G1468gat, G1370gat);
nand NAND2_280 (G1469gat, G1370gat, G1222gat);
not NOT1_281 (G1470gat, G1376gat);
nand NAND2_282 (G1471gat, G1376gat, G1227gat);
nand NAND2_283 (G1472gat, G1387gat, G1433gat);
not NOT1_284 (G1475gat, G1390gat);
nand NAND2_285 (G1476gat, G1390gat, G1240gat);
nand NAND2_286 (G1478gat, G1389gat, G1434gat);
nand NAND2_287 (G1481gat, G1399gat, G1439gat);
nand NAND2_288 (G1484gat, G1397gat, G1438gat);
nand NAND2_289 (G1487gat, G939gat, G1444gat);
nand NAND2_290 (G1488gat, G935gat, G1446gat);
nand NAND2_291 (G1489gat, G943gat, G1448gat);
not NOT1_292 (G1490gat, G1419gat);
not NOT1_293 (G1491gat, G1416gat);
nand NAND2_294 (G1492gat, G947gat, G1452gat);
nand NAND2_295 (G1493gat, G955gat, G1454gat);
nand NAND2_296 (G1494gat, G951gat, G1456gat);
nand NAND2_297 (G1495gat, G969gat, G1458gat);
nand NAND2_298 (G1496gat, G977gat, G1460gat);
nand NAND2_299 (G1498gat, G998gat, G1463gat);
not NOT1_300 (G1499gat, G1440gat);
nand NAND2_301 (G1500gat, G965gat, G1468gat);
nand NAND2_302 (G1501gat, G973gat, G1470gat);
nand NAND2_303 (G1504gat, G994gat, G1475gat);
not NOT1_304 (G1510gat, G1464gat);
nand NAND2_305 (G1513gat, G1443gat, G1487gat);
nand NAND2_306 (G1514gat, G1445gat, G1488gat);
nand NAND2_307 (G1517gat, G1447gat, G1489gat);
nand NAND2_308 (G1520gat, G1451gat, G1492gat);
nand NAND2_309 (G1521gat, G1453gat, G1493gat);
nand NAND2_310 (G1522gat, G1455gat, G1494gat);
nand NAND2_311 (G1526gat, G1457gat, G1495gat);
nand NAND2_312 (G1527gat, G1459gat, G1496gat);
not NOT1_313 (G1528gat, G1472gat);
nand NAND2_314 (G1529gat, G1462gat, G1498gat);
not NOT1_315 (G1530gat, G1478gat);
not NOT1_316 (G1531gat, G1481gat);
not NOT1_317 (G1532gat, G1484gat);
nand NAND2_318 (G1534gat, G1471gat, G1501gat);
nand NAND2_319 (G1537gat, G1469gat, G1500gat);
nand NAND2_320 (G1540gat, G1476gat, G1504gat);
not NOT1_321 (G1546gat, G1513gat);
not NOT1_322 (G1554gat, G1521gat);
not NOT1_323 (G1557gat, G1526gat);
not NOT1_324 (G1561gat, G1520gat);
nand NAND2_325 (G1567gat, G1484gat, G1531gat);
nand NAND2_326 (G1568gat, G1481gat, G1532gat);
not NOT1_327 (G1569gat, G1510gat);
not NOT1_328 (G1571gat, G1527gat);
not NOT1_329 (G1576gat, G1529gat);
not NOT1_330 (G1591gat, G1534gat);
not NOT1_331 (G1593gat, G1537gat);
nand NAND2_332 (G1594gat, G1540gat, G1530gat);
not NOT1_333 (G1595gat, G1540gat);
nand NAND2_334 (G1596gat, G1567gat, G1568gat);
not NOT1_335 (G1635gat, G1571gat);
nand NAND2_336 (G1636gat, G1478gat, G1595gat);
nand NAND2_337 (G1638gat, G1576gat, G1569gat);
not NOT1_338 (G1639gat, G1576gat);
nand NAND2_339 (G1671gat, G1596gat, G893gat);
not NOT1_340 (G1672gat, G1596gat);
not NOT1_341 (G1675gat, G1600gat);
not NOT1_342 (G1677gat, G1603gat);
nand NAND2_343 (G1678gat, G1606gat, G1217gat);
not NOT1_344 (G1679gat, G1606gat);
nand NAND2_345 (G1680gat, G1609gat, G1219gat);
not NOT1_346 (G1681gat, G1609gat);
not NOT1_347 (G1682gat, G1612gat);
not NOT1_348 (G1683gat, G1615gat);
nand NAND2_349 (G1685gat, G1594gat, G1636gat);
nand NAND2_350 (G1688gat, G1510gat, G1639gat);
nand NAND2_351 (G1706gat, G643gat, G1672gat);
not NOT1_352 (G1707gat, G1643gat);
nand NAND2_353 (G1708gat, G1647gat, G1675gat);
not NOT1_354 (G1709gat, G1647gat);
nand NAND2_355 (G1710gat, G1651gat, G1677gat);
not NOT1_356 (G1711gat, G1651gat);
nand NAND2_357 (G1712gat, G1028gat, G1679gat);
nand NAND2_358 (G1713gat, G1031gat, G1681gat);
nand NAND2_359 (G1720gat, G1658gat, G1593gat);
not NOT1_360 (G1721gat, G1658gat);
nand NAND2_361 (G1723gat, G1638gat, G1688gat);
not NOT1_362 (G1727gat, G1661gat);
not NOT1_363 (G1728gat, G1640gat);
not NOT1_364 (G1730gat, G1664gat);
nand NAND2_365 (G1740gat, G1685gat, G1528gat);
not NOT1_366 (G1741gat, G1685gat);
nand NAND2_367 (G1742gat, G1671gat, G1706gat);
nand NAND2_368 (G1746gat, G1600gat, G1709gat);
nand NAND2_369 (G1747gat, G1603gat, G1711gat);
nand NAND2_370 (G1748gat, G1678gat, G1712gat);
nand NAND2_371 (G1751gat, G1680gat, G1713gat);
nand NAND2_372 (G1759gat, G1537gat, G1721gat);
not NOT1_373 (G1761gat, G1697gat);
nand NAND2_374 (G1762gat, G1697gat, G1727gat);
not NOT1_375 (G1763gat, G1701gat);
nand NAND2_376 (G1764gat, G1701gat, G1730gat);
not NOT1_377 (G1768gat, G1717gat);
nand NAND2_378 (G1769gat, G1472gat, G1741gat);
nand NAND2_379 (G1772gat, G1723gat, G1413gat);
not NOT1_380 (G1773gat, G1723gat);
nand NAND2_381 (G1774gat, G1708gat, G1746gat);
nand NAND2_382 (G1777gat, G1710gat, G1747gat);
not NOT1_383 (G1783gat, G1731gat);
nand NAND2_384 (G1784gat, G1731gat, G1682gat);
not NOT1_385 (G1785gat, G1714gat);
not NOT1_386 (G1786gat, G1734gat);
nand NAND2_387 (G1787gat, G1734gat, G1683gat);
nand NAND2_388 (G1788gat, G1720gat, G1759gat);
nand NAND2_389 (G1791gat, G1661gat, G1761gat);
nand NAND2_390 (G1792gat, G1664gat, G1763gat);
nand NAND2_391 (G1795gat, G1751gat, G1155gat);
not NOT1_392 (G1796gat, G1751gat);
nand NAND2_393 (G1798gat, G1740gat, G1769gat);
nand NAND2_394 (G1801gat, G1334gat, G1773gat);
nand NAND2_395 (G1802gat, G1742gat, G290gat);
not NOT1_396 (G1807gat, G1748gat);
nand NAND2_397 (G1808gat, G1748gat, G1218gat);
nand NAND2_398 (G1809gat, G1612gat, G1783gat);
nand NAND2_399 (G1810gat, G1615gat, G1786gat);
nand NAND2_400 (G1812gat, G1791gat, G1762gat);
nand NAND2_401 (G1815gat, G1792gat, G1764gat);
nand NAND2_402 (G1821gat, G1777gat, G1490gat);
not NOT1_403 (G1822gat, G1777gat);
nand NAND2_404 (G1823gat, G1774gat, G1491gat);
not NOT1_405 (G1824gat, G1774gat);
nand NAND2_406 (G1825gat, G962gat, G1796gat);
nand NAND2_407 (G1826gat, G1788gat, G1409gat);
not NOT1_408 (G1827gat, G1788gat);
nand NAND2_409 (G1830gat, G1772gat, G1801gat);
nand NAND2_410 (G1837gat, G959gat, G1807gat);
nand NAND2_411 (G1838gat, G1809gat, G1784gat);
nand NAND2_412 (G1841gat, G1810gat, G1787gat);
nand NAND2_413 (G1848gat, G1419gat, G1822gat);
nand NAND2_414 (G1849gat, G1416gat, G1824gat);
nand NAND2_415 (G1850gat, G1795gat, G1825gat);
nand NAND2_416 (G1852gat, G1319gat, G1827gat);
nand NAND2_417 (G1855gat, G1815gat, G1707gat);
not NOT1_418 (G1856gat, G1815gat);
not NOT1_419 (G1857gat, G1818gat);
nand NAND2_420 (G1858gat, G1798gat, G290gat);
not NOT1_421 (G1864gat, G1812gat);
nand NAND2_422 (G1865gat, G1812gat, G1728gat);
nand NAND2_423 (G1875gat, G1808gat, G1837gat);
nand NAND2_424 (G1878gat, G1821gat, G1848gat);
nand NAND2_425 (G1879gat, G1823gat, G1849gat);
nand NAND2_426 (G1882gat, G1841gat, G1768gat);
not NOT1_427 (G1883gat, G1841gat);
nand NAND2_428 (G1884gat, G1826gat, G1852gat);
nand NAND2_429 (G1885gat, G1643gat, G1856gat);
nand NAND2_430 (G1889gat, G1830gat, G290gat);
not NOT1_431 (G1895gat, G1838gat);
nand NAND2_432 (G1896gat, G1838gat, G1785gat);
nand NAND2_433 (G1897gat, G1640gat, G1864gat);
not NOT1_434 (G1898gat, G1850gat);
not NOT1_435 (G1910gat, G1878gat);
nand NAND2_436 (G1911gat, G1717gat, G1883gat);
not NOT1_437 (G1912gat, G1884gat);
nand NAND2_438 (G1913gat, G1855gat, G1885gat);
not NOT1_439 (G1915gat, G1866gat);
nand NAND2_440 (G1919gat, G1872gat, G919gat);
not NOT1_441 (G1920gat, G1872gat);
nand NAND2_442 (G1921gat, G1869gat, G920gat);
not NOT1_443 (G1922gat, G1869gat);
not NOT1_444 (G1923gat, G1875gat);
nand NAND2_445 (G1924gat, G1714gat, G1895gat);
nand NAND2_446 (G1933gat, G1865gat, G1897gat);
nand NAND2_447 (G1936gat, G1882gat, G1911gat);
not NOT1_448 (G1937gat, G1898gat);
not NOT1_449 (G1938gat, G1902gat);
nand NAND2_450 (G1941gat, G679gat, G1920gat);
nand NAND2_451 (G1942gat, G676gat, G1922gat);
not NOT1_452 (G1947gat, G1913gat);
nand NAND2_453 (G1961gat, G1896gat, G1924gat);
and AND2_454 (G1965gat, G1910gat, G601gat);
and AND2_455 (G1968gat, G602gat, G1912gat);
nand NAND2_456 (G1975gat, G1930gat, G917gat);
not NOT1_457 (G1976gat, G1930gat);
nand NAND2_458 (G1977gat, G1927gat, G918gat);
not NOT1_459 (G1978gat, G1927gat);
nand NAND2_460 (G1979gat, G1919gat, G1941gat);
nand NAND2_461 (G1980gat, G1921gat, G1942gat);
not NOT1_462 (G1985gat, G1933gat);
not NOT1_463 (G1987gat, G1936gat);
not NOT1_464 (G1999gat, G1944gat);
nand NAND2_465 (G2000gat, G1944gat, G1937gat);
not NOT1_466 (G2002gat, G1947gat);
nand NAND2_467 (G2003gat, G1947gat, G1499gat);
nand NAND2_468 (G2004gat, G1953gat, G1350gat);
not NOT1_469 (G2005gat, G1953gat);
nand NAND2_470 (G2006gat, G1950gat, G1351gat);
not NOT1_471 (G2007gat, G1950gat);
nand NAND2_472 (G2008gat, G673gat, G1976gat);
nand NAND2_473 (G2009gat, G670gat, G1978gat);
not NOT1_474 (G2012gat, G1979gat);
not NOT1_475 (G2013gat, G1958gat);
nand NAND2_476 (G2014gat, G1958gat, G1923gat);
not NOT1_477 (G2015gat, G1961gat);
nand NAND2_478 (G2016gat, G1961gat, G1635gat);
not NOT1_479 (G2018gat, G1965gat);
not NOT1_480 (G2019gat, G1968gat);
nand NAND2_481 (G2020gat, G1898gat, G1999gat);
not NOT1_482 (G2021gat, G1987gat);
nand NAND2_483 (G2022gat, G1987gat, G1591gat);
nand NAND2_484 (G2023gat, G1440gat, G2002gat);
nand NAND2_485 (G2024gat, G1261gat, G2005gat);
nand NAND2_486 (G2025gat, G1258gat, G2007gat);
nand NAND2_487 (G2026gat, G1975gat, G2008gat);
nand NAND2_488 (G2027gat, G1977gat, G2009gat);
not NOT1_489 (G2030gat, G1980gat);
nand NAND2_490 (G2036gat, G1875gat, G2013gat);
nand NAND2_491 (G2037gat, G1571gat, G2015gat);
nand NAND2_492 (G2038gat, G2020gat, G2000gat);
nand NAND2_493 (G2039gat, G1534gat, G2021gat);
nand NAND2_494 (G2040gat, G2023gat, G2003gat);
nand NAND2_495 (G2041gat, G2004gat, G2024gat);
nand NAND2_496 (G2042gat, G2006gat, G2025gat);
not NOT1_497 (G2047gat, G2026gat);
nand NAND2_498 (G2052gat, G2036gat, G2014gat);
nand NAND2_499 (G2055gat, G2037gat, G2016gat);
not NOT1_500 (G2060gat, G2038gat);
nand NAND2_501 (G2061gat, G2039gat, G2022gat);
nand NAND2_502 (G2062gat, G2040gat, G290gat);
not NOT1_503 (G2067gat, G2041gat);
not NOT1_504 (G2068gat, G2027gat);
not NOT1_505 (G2076gat, G2052gat);
not NOT1_506 (G2077gat, G2055gat);
nand NAND2_507 (G2078gat, G2060gat, G290gat);
nand NAND2_508 (G2081gat, G2061gat, G290gat);
not NOT1_509 (G2086gat, G2042gat);
and AND2_510 (G2104gat, G2030gat, G2068gat);
and AND2_511 (G2119gat, G2033gat, G2068gat);
and AND2_512 (G2129gat, G2030gat, G2071gat);
and AND2_513 (G2143gat, G2033gat, G2071gat);
nand NAND2_514 (G2214gat, G2151gat, G915gat);
not NOT1_515 (G2215gat, G2151gat);
nand NAND2_516 (G2216gat, G2148gat, G916gat);
not NOT1_517 (G2217gat, G2148gat);
nand NAND2_518 (G2222gat, G2199gat, G1348gat);
not NOT1_519 (G2223gat, G2199gat);
nand NAND2_520 (G2224gat, G2196gat, G1349gat);
not NOT1_521 (G2225gat, G2196gat);
nand NAND2_522 (G2226gat, G2205gat, G913gat);
not NOT1_523 (G2227gat, G2205gat);
nand NAND2_524 (G2228gat, G2202gat, G914gat);
not NOT1_525 (G2229gat, G2202gat);
nand NAND2_526 (G2230gat, G667gat, G2215gat);
nand NAND2_527 (G2231gat, G664gat, G2217gat);
nand NAND2_528 (G2232gat, G1255gat, G2223gat);
nand NAND2_529 (G2233gat, G1252gat, G2225gat);
nand NAND2_530 (G2234gat, G661gat, G2227gat);
nand NAND2_531 (G2235gat, G658gat, G2229gat);
nand NAND2_532 (G2236gat, G2214gat, G2230gat);
nand NAND2_533 (G2237gat, G2216gat, G2231gat);
nand NAND2_534 (G2240gat, G2222gat, G2232gat);
nand NAND2_535 (G2241gat, G2224gat, G2233gat);
nand NAND2_536 (G2244gat, G2226gat, G2234gat);
nand NAND2_537 (G2245gat, G2228gat, G2235gat);
not NOT1_538 (G2250gat, G2236gat);
not NOT1_539 (G2253gat, G2240gat);
not NOT1_540 (G2256gat, G2244gat);
not NOT1_541 (G2257gat, G2237gat);
not NOT1_542 (G2263gat, G2241gat);
and AND2_543 (G2266gat, G1164gat, G2241gat);
not NOT1_544 (G2269gat, G2245gat);
and AND2_545 (G2272gat, G1168gat, G2245gat);
and AND4_546 (G2273gat, G2067gat, G2012gat, G2047gat, G2250gat);
and AND4_547 (G2274gat, G899gat, G2256gat, G2253gat, G903gat);
nand NAND2_548 (G2279gat, G2273gat, G2274gat);
and AND2_549 (G2340gat, G2086gat, G2257gat);
and AND2_550 (G2353gat, G2089gat, G2257gat);
and AND2_551 (G2361gat, G2086gat, G2260gat);
and AND2_552 (G2375gat, G2089gat, G2260gat);
and AND4_553 (G2384gat, G338gat, G2279gat, G313gat, G313gat);
and AND2_554 (G2385gat, G1163gat, G2263gat);
and AND2_555 (G2386gat, G1164gat, G2263gat);
and AND2_556 (G2426gat, G1167gat, G2269gat);
and AND2_557 (G2427gat, G1168gat, G2269gat);
nand NAND5_558 (G2537gat, G2286gat, G2315gat, G2361gat, G2104gat, G1171gat);
nand NAND5_559 (G2540gat, G2286gat, G2315gat, G2340gat, G2129gat, G1171gat);
nand NAND5_560 (G2543gat, G2286gat, G2315gat, G2340gat, G2119gat, G1171gat);
nand NAND5_561 (G2546gat, G2286gat, G2315gat, G2353gat, G2104gat, G1171gat);
nand NAND5_562 (G2549gat, G2297gat, G2315gat, G2375gat, G2119gat, G1188gat);
nand NAND5_563 (G2552gat, G2297gat, G2326gat, G2361gat, G2143gat, G1188gat);
nand NAND5_564 (G2555gat, G2297gat, G2326gat, G2375gat, G2129gat, G1188gat);
and AND5_565 (G2558gat, G2286gat, G2315gat, G2361gat, G2104gat, G1171gat);
and AND5_566 (G2561gat, G2286gat, G2315gat, G2340gat, G2129gat, G1171gat);
and AND5_567 (G2564gat, G2286gat, G2315gat, G2340gat, G2119gat, G1171gat);
and AND5_568 (G2567gat, G2286gat, G2315gat, G2353gat, G2104gat, G1171gat);
and AND5_569 (G2570gat, G2297gat, G2315gat, G2375gat, G2119gat, G1188gat);
and AND5_570 (G2573gat, G2297gat, G2326gat, G2361gat, G2143gat, G1188gat);
and AND5_571 (G2576gat, G2297gat, G2326gat, G2375gat, G2129gat, G1188gat);
nand NAND5_572 (G2594gat, G2286gat, G2427gat, G2361gat, G2129gat, G1171gat);
nand NAND5_573 (G2597gat, G2297gat, G2427gat, G2361gat, G2119gat, G1171gat);
nand NAND5_574 (G2600gat, G2297gat, G2427gat, G2375gat, G2104gat, G1171gat);
nand NAND5_575 (G2603gat, G2297gat, G2427gat, G2340gat, G2143gat, G1171gat);
nand NAND5_576 (G2606gat, G2297gat, G2427gat, G2353gat, G2129gat, G1188gat);
nand NAND5_577 (G2611gat, G2386gat, G2326gat, G2361gat, G2129gat, G1188gat);
nand NAND5_578 (G2614gat, G2386gat, G2326gat, G2361gat, G2119gat, G1188gat);
nand NAND5_579 (G2617gat, G2386gat, G2326gat, G2375gat, G2104gat, G1188gat);
nand NAND5_580 (G2620gat, G2386gat, G2326gat, G2353gat, G2129gat, G1188gat);
nand NAND5_581 (G2627gat, G2297gat, G2427gat, G2340gat, G2104gat, G926gat);
nand NAND5_582 (G2628gat, G2386gat, G2326gat, G2340gat, G2104gat, G926gat);
nand NAND5_583 (G2629gat, G2386gat, G2427gat, G2361gat, G2104gat, G926gat);
nand NAND5_584 (G2630gat, G2386gat, G2427gat, G2340gat, G2129gat, G926gat);
nand NAND5_585 (G2631gat, G2386gat, G2427gat, G2340gat, G2119gat, G926gat);
nand NAND5_586 (G2632gat, G2386gat, G2427gat, G2353gat, G2104gat, G926gat);
nand NAND5_587 (G2633gat, G2386gat, G2426gat, G2340gat, G2104gat, G926gat);
nand NAND5_588 (G2634gat, G2385gat, G2427gat, G2340gat, G2104gat, G926gat);
and AND5_589 (G2639gat, G2286gat, G2427gat, G2361gat, G2129gat, G1171gat);
and AND5_590 (G2642gat, G2297gat, G2427gat, G2361gat, G2119gat, G1171gat);
and AND5_591 (G2645gat, G2297gat, G2427gat, G2375gat, G2104gat, G1171gat);
and AND5_592 (G2648gat, G2297gat, G2427gat, G2340gat, G2143gat, G1171gat);
and AND5_593 (G2651gat, G2297gat, G2427gat, G2353gat, G2129gat, G1188gat);
and AND5_594 (G2655gat, G2386gat, G2326gat, G2361gat, G2129gat, G1188gat);
and AND5_595 (G2658gat, G2386gat, G2326gat, G2361gat, G2119gat, G1188gat);
and AND5_596 (G2661gat, G2386gat, G2326gat, G2375gat, G2104gat, G1188gat);
and AND5_597 (G2664gat, G2386gat, G2326gat, G2353gat, G2129gat, G1188gat);
nand NAND2_598 (G2669gat, G2558gat, G534gat);
not NOT1_599 (G2670gat, G2558gat);
nand NAND2_600 (G2671gat, G2561gat, G535gat);
not NOT1_601 (G2672gat, G2561gat);
nand NAND2_602 (G2673gat, G2564gat, G536gat);
not NOT1_603 (G2674gat, G2564gat);
nand NAND2_604 (G2675gat, G2567gat, G537gat);
not NOT1_605 (G2676gat, G2567gat);
nand NAND2_606 (G2682gat, G2570gat, G543gat);
not NOT1_607 (G2683gat, G2570gat);
nand NAND2_608 (G2688gat, G2573gat, G548gat);
not NOT1_609 (G2689gat, G2573gat);
nand NAND2_610 (G2690gat, G2576gat, G549gat);
not NOT1_611 (G2691gat, G2576gat);
and AND4_612 (G2692gat, G2627gat, G2628gat, G2629gat, G2630gat);
and AND4_613 (G2693gat, G2631gat, G2632gat, G2633gat, G2634gat);
and AND2_614 (G2710gat, G2692gat, G2693gat);
nand NAND2_615 (G2720gat, G343gat, G2670gat);
nand NAND2_616 (G2721gat, G346gat, G2672gat);
nand NAND2_617 (G2722gat, G349gat, G2674gat);
nand NAND2_618 (G2723gat, G352gat, G2676gat);
nand NAND2_619 (G2724gat, G2639gat, G538gat);
not NOT1_620 (G2725gat, G2639gat);
nand NAND2_621 (G2726gat, G2642gat, G539gat);
not NOT1_622 (G2727gat, G2642gat);
nand NAND2_623 (G2728gat, G2645gat, G540gat);
not NOT1_624 (G2729gat, G2645gat);
nand NAND2_625 (G2730gat, G2648gat, G541gat);
not NOT1_626 (G2731gat, G2648gat);
nand NAND2_627 (G2732gat, G2651gat, G542gat);
not NOT1_628 (G2733gat, G2651gat);
nand NAND2_629 (G2734gat, G370gat, G2683gat);
nand NAND2_630 (G2735gat, G2655gat, G544gat);
not NOT1_631 (G2736gat, G2655gat);
nand NAND2_632 (G2737gat, G2658gat, G545gat);
not NOT1_633 (G2738gat, G2658gat);
nand NAND2_634 (G2739gat, G2661gat, G546gat);
not NOT1_635 (G2740gat, G2661gat);
nand NAND2_636 (G2741gat, G2664gat, G547gat);
not NOT1_637 (G2742gat, G2664gat);
nand NAND2_638 (G2743gat, G385gat, G2689gat);
nand NAND2_639 (G2744gat, G388gat, G2691gat);
and AND4_640 (G27440gat, G2537gat, G2540gat, G2543gat, G2546gat);
and AND4_641 (G27441gat, G2594gat, G2597gat, G2600gat, G2603gat);
nand NAND2_642 (G2745gat, G27440gat, G27441gat);
and AND4_643 (G27450gat, G2606gat, G2549gat, G2611gat, G2614gat);
and AND4_644 (G27451gat, G2617gat, G2620gat, G2552gat, G2555gat);
nand NAND2_645 (G2746gat, G27450gat, G27451gat);
and AND4_646 (G27460gat, G2537gat, G2540gat, G2543gat, G2546gat);
and AND4_647 (G27461gat, G2594gat, G2597gat, G2600gat, G2603gat);
and AND2_648 (G2747gat, G27460gat, G27461gat);
and AND4_649 (G27470gat, G2606gat, G2549gat, G2611gat, G2614gat);
and AND4_650 (G27471gat, G2617gat, G2620gat, G2552gat, G2555gat);
and AND2_651 (G2750gat, G27470gat, G27471gat);
nand NAND2_652 (G2753gat, G2669gat, G2720gat);
nand NAND2_653 (G2754gat, G2671gat, G2721gat);
nand NAND2_654 (G2755gat, G2673gat, G2722gat);
nand NAND2_655 (G2756gat, G2675gat, G2723gat);
nand NAND2_656 (G2757gat, G355gat, G2725gat);
nand NAND2_657 (G2758gat, G358gat, G2727gat);
nand NAND2_658 (G2759gat, G361gat, G2729gat);
nand NAND2_659 (G2760gat, G364gat, G2731gat);
nand NAND2_660 (G2761gat, G367gat, G2733gat);
nand NAND2_661 (G2762gat, G2682gat, G2734gat);
nand NAND2_662 (G2763gat, G373gat, G2736gat);
nand NAND2_663 (G2764gat, G376gat, G2738gat);
nand NAND2_664 (G2765gat, G379gat, G2740gat);
nand NAND2_665 (G2766gat, G382gat, G2742gat);
nand NAND2_666 (G2767gat, G2688gat, G2743gat);
nand NAND2_667 (G2768gat, G2690gat, G2744gat);
and AND2_668 (G2773gat, G2745gat, G275gat);
and AND2_669 (G2776gat, G2746gat, G276gat);
nand NAND2_670 (G2779gat, G2724gat, G2757gat);
nand NAND2_671 (G2780gat, G2726gat, G2758gat);
nand NAND2_672 (G2781gat, G2728gat, G2759gat);
nand NAND2_673 (G2782gat, G2730gat, G2760gat);
nand NAND2_674 (G2783gat, G2732gat, G2761gat);
nand NAND2_675 (G2784gat, G2735gat, G2763gat);
nand NAND2_676 (G2785gat, G2737gat, G2764gat);
nand NAND2_677 (G2786gat, G2739gat, G2765gat);
nand NAND2_678 (G2787gat, G2741gat, G2766gat);
and AND3_679 (G2788gat, G2747gat, G2750gat, G2710gat);
nand NAND2_680 (G2789gat, G2747gat, G2750gat);
and AND4_681 (G2800gat, G338gat, G2279gat, G99gat, G2788gat);
nand NAND2_682 (G2807gat, G2773gat, G2018gat);
not NOT1_683 (G2808gat, G2773gat);
nand NAND2_684 (G2809gat, G2776gat, G2019gat);
not NOT1_685 (G2810gat, G2776gat);
nor NOR2_686 (G2811gat, G2384gat, G2800gat);
and AND3_687 (G2812gat, G897gat, G283gat, G2789gat);
and AND3_688 (G2815gat, G76gat, G283gat, G2789gat);
and AND3_689 (G2818gat, G82gat, G283gat, G2789gat);
and AND3_690 (G2821gat, G85gat, G283gat, G2789gat);
and AND3_691 (G2824gat, G898gat, G283gat, G2789gat);
nand NAND2_692 (G2827gat, G1965gat, G2808gat);
nand NAND2_693 (G2828gat, G1968gat, G2810gat);
and AND3_694 (G2829gat, G79gat, G283gat, G2789gat);
nand NAND2_695 (G2843gat, G2807gat, G2827gat);
nand NAND2_696 (G2846gat, G2809gat, G2828gat);
nand NAND2_697 (G2850gat, G2812gat, G2076gat);
nand NAND2_698 (G2851gat, G2815gat, G2077gat);
nand NAND2_699 (G2852gat, G2818gat, G1915gat);
nand NAND2_700 (G2853gat, G2821gat, G1857gat);
nand NAND2_701 (G2854gat, G2824gat, G1938gat);
not NOT1_702 (G2857gat, G2812gat);
not NOT1_703 (G2858gat, G2815gat);
not NOT1_704 (G2859gat, G2818gat);
not NOT1_705 (G2860gat, G2821gat);
not NOT1_706 (G2861gat, G2824gat);
not NOT1_707 (G2862gat, G2829gat);
nand NAND2_708 (G2863gat, G2829gat, G1985gat);
nand NAND2_709 (G2866gat, G2052gat, G2857gat);
nand NAND2_710 (G2867gat, G2055gat, G2858gat);
nand NAND2_711 (G2868gat, G1866gat, G2859gat);
nand NAND2_712 (G2869gat, G1818gat, G2860gat);
nand NAND2_713 (G2870gat, G1902gat, G2861gat);
nand NAND2_714 (G2871gat, G2843gat, G886gat);
not NOT1_715 (G2872gat, G2843gat);
nand NAND2_716 (G2873gat, G2846gat, G887gat);
not NOT1_717 (G2874gat, G2846gat);
nand NAND2_718 (G2875gat, G1933gat, G2862gat);
nand NAND2_719 (G2876gat, G2866gat, G2850gat);
nand NAND2_720 (G2877gat, G2867gat, G2851gat);
nand NAND2_721 (G2878gat, G2868gat, G2852gat);
nand NAND2_722 (G2879gat, G2869gat, G2853gat);
nand NAND2_723 (G2880gat, G2870gat, G2854gat);
nand NAND2_724 (G2881gat, G682gat, G2872gat);
nand NAND2_725 (G2882gat, G685gat, G2874gat);
nand NAND2_726 (G2883gat, G2875gat, G2863gat);
and AND2_727 (G2886gat, G2876gat, G550gat);
and AND2_728 (G2887gat, G551gat, G2877gat);
and AND2_729 (G2888gat, G553gat, G2878gat);
and AND2_730 (G2889gat, G2879gat, G554gat);
and AND2_731 (G2890gat, G555gat, G2880gat);
nand NAND2_732 (G2891gat, G2871gat, G2881gat);
nand NAND2_733 (G2892gat, G2873gat, G2882gat);
nand NAND2_734 (G2895gat, G2883gat, G1461gat);
not NOT1_735 (G2896gat, G2883gat);
nand NAND2_736 (G2897gat, G1383gat, G2896gat);
nand NAND2_737 (G2898gat, G2895gat, G2897gat);
and AND2_738 (G2899gat, G2898gat, G552gat);

endmodule