module c3540_sarlock_8k(G1gat,G13gat,G20gat,G33gat,G41gat,G45gat,G50gat,G58gat,G68gat,G77gat,G87gat,G97gat,G107gat,G116gat,G124gat,G125gat,G128gat,G132gat,G137gat,G143gat,G150gat,G159gat,G169gat,G179gat,G190gat,G200gat,G213gat,G222gat,G223gat,G226gat,G232gat,G238gat,G244gat,G250gat,G257gat,G264gat,G270gat,G274gat,G283gat,G294gat,G303gat,G311gat,G317gat,G322gat,G326gat,G329gat,G330gat,G343gat,G349gat,G350gat,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,G1713gat,G1947gat,G3195gat,G3833gat,G3987gat,G4028gat,G4145gat,G4589gat,G4667gat,G4815gat,G4944gat,G5002gat,G5045gat,G5047gat,G5078gat,G5102gat,G5120gat,G5121gat,G5192gat,G5231gat,G5360gat,G5361gat);

input G1gat,G13gat,G20gat,G33gat,G41gat,G45gat,G50gat,G58gat,G68gat,G77gat,G87gat,G97gat,G107gat,G116gat,G124gat,G125gat,G128gat,G132gat,G137gat,G143gat,G150gat,G159gat,G169gat,G179gat,G190gat,G200gat,G213gat,G222gat,G223gat,G226gat,G232gat,G238gat,G244gat,G250gat,G257gat,G264gat,G270gat,G274gat,G283gat,G294gat,G303gat,G311gat,G317gat,G322gat,G326gat,G329gat,G330gat,G343gat,G349gat,G350gat,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7;
output G1713gat,G1947gat,G3195gat,G3833gat,G3987gat,G4028gat,G4145gat,G4589gat,G4667gat,G4815gat,G4944gat,G5002gat,G5045gat,G5047gat,G5078gat,G5102gat,G5120gat,G5121gat,G5192gat,G5231gat,G5360gat,G5361gat;
wire G665gat,G679gat,G686gat,G702gat,G724gat,G736gat,G749gat,G763gat,G768gat,G769gat,G779gat,G786gat,G793gat,G794gat,G803gat,G820gat,G825gat,G829gat,G832gat,G835gat,G839gat,G842gat,G848gat,G854gat,G861gat,G867gat,G870gat,G883gat,G889gat,G890gat,G891gat,G892gat,G895gat,G896gat,G913gat,G914gat,G915gat,G916gat,G920gat,G1067gat,G1117gat,G1179gat,G1196gat,G1197gat,G1202gat,G1219gat,G1250gat,G1251gat,G1252gat,G1253gat,G1254gat,G1255gat,G1256gat,G1257gat,G1258gat,G1259gat,G1260gat,G1261gat,G1262gat,G1263gat,G1264gat,G1267gat,G1271gat,G1272gat,G1306gat,G1315gat,G1322gat,G1325gat,G1328gat,G1331gat,G1337gat,G1338gat,G1339gat,G1340gat,G1343gat,G1344gat,G1345gat,G1346gat,G1347gat,G1348gat,G1349gat,G1350gat,G1351gat,G1352gat,G1353gat,G1358gat,G1366gat,G1401gat,G1402gat,G1403gat,G1404gat,G1405gat,G1406gat,G1407gat,G1408gat,G1409gat,G1426gat,G1427gat,G1452gat,G1459gat,G1460gat,G1461gat,G1464gat,G1467gat,G1468gat,G1469gat,G1470gat,G1474gat,G1505gat,G1507gat,G1508gat,G1509gat,G1510gat,G1511gat,G1512gat,G1520gat,G1562gat,G1579gat,G1580gat,G1581gat,G1582gat,G1583gat,G1584gat,G1585gat,G1586gat,G1587gat,G1588gat,G1589gat,G1590gat,G1591gat,G1592gat,G1593gat,G1594gat,G1595gat,G1596gat,G1597gat,G1598gat,G1599gat,G1600gat,G1643gat,G1644gat,G1645gat,G1646gat,G1647gat,G1648gat,G1649gat,G1650gat,G1667gat,G1670gat,G1673gat,G1674gat,G1675gat,G1676gat,G1677gat,G1678gat,G1679gat,G1680gat,G1691gat,G1692gat,G1693gat,G1694gat,G1714gat,G1715gat,G1718gat,G1721gat,G1722gat,G1725gat,G1726gat,G1727gat,G1728gat,G1729gat,G1730gat,G1731gat,G1735gat,G1736gat,G1737gat,G1738gat,G1747gat,G1756gat,G1761gat,G1764gat,G1765gat,G1766gat,G1767gat,G1768gat,G1769gat,G1770gat,G1787gat,G1788gat,G1789gat,G1790gat,G1791gat,G1792gat,G1793gat,G1794gat,G1795gat,G1796gat,G1797gat,G1798gat,G1799gat,G1800gat,G1801gat,G1802gat,G1803gat,G1806gat,G1809gat,G1812gat,G1815gat,G1818gat,G1821gat,G1824gat,G1833gat,G1842gat,G1843gat,G1844gat,G1845gat,G1846gat,G1847gat,G1848gat,G1849gat,G1850gat,G1851gat,G1852gat,G1853gat,G1854gat,G1855gat,G1856gat,G1857gat,G1858gat,G1859gat,G1860gat,G1861gat,G1862gat,G1863gat,G1864gat,G1869gat,G1870gat,G1873gat,G1874gat,G1875gat,G1878gat,G1879gat,G1880gat,G1883gat,G1884gat,G1885gat,G1888gat,G1889gat,G1890gat,G1893gat,G1894gat,G1895gat,G1898gat,G1899gat,G1900gat,G1903gat,G1904gat,G1905gat,G1908gat,G1909gat,G1912gat,G1913gat,G1917gat,G1922gat,G1926gat,G1933gat,G1936gat,G1939gat,G1940gat,G1941gat,G1942gat,G1943gat,G1944gat,G1945gat,G1946gat,G1960gat,G1961gat,G1966gat,G1981gat,G1982gat,G1983gat,G1986gat,G1987gat,G1988gat,G1989gat,G1990gat,G1991gat,G2022gat,G2023gat,G2024gat,G2025gat,G2026gat,G2027gat,G2028gat,G2029gat,G2030gat,G2031gat,G2032gat,G2033gat,G2034gat,G2035gat,G2036gat,G2037gat,G2043gat,G2057gat,G2068gat,G2073gat,G2078gat,G2083gat,G2088gat,G2093gat,G2098gat,G2103gat,G2121gat,G2122gat,G2123gat,G2124gat,G2125gat,G2126gat,G2127gat,G2128gat,G2133gat,G2134gat,G2135gat,G2136gat,G2137gat,G2138gat,G2139gat,G2141gat,G2142gat,G2143gat,G2144gat,G2145gat,G2146gat,G2147gat,G2148gat,G2149gat,G2150gat,G2151gat,G2152gat,G2153gat,G2154gat,G2155gat,G2156gat,G2157gat,G2178gat,G2179gat,G2180gat,G2181gat,G2183gat,G2184gat,G2185gat,G2188gat,G2191gat,G2194gat,G2197gat,G2200gat,G2203gat,G2206gat,G2209gat,G2210gat,G2211gat,G2230gat,G2231gat,G2232gat,G2233gat,G2234gat,G2235gat,G2236gat,G2237gat,G2238gat,G2239gat,G2240gat,G2241gat,G2242gat,G2243gat,G2244gat,G2245gat,G2270gat,G2277gat,G2282gat,G2287gat,G2294gat,G2299gat,G2307gat,G2310gat,G2325gat,G2328gat,G2331gat,G2334gat,G2341gat,G2342gat,G2347gat,G2348gat,G2349gat,G2350gat,G2351gat,G2352gat,G2353gat,G2354gat,G2355gat,G2374gat,G2375gat,G2376gat,G2379gat,G2398gat,G2417gat,G2418gat,G2419gat,G2420gat,G2421gat,G2422gat,G2425gat,G2426gat,G2427gat,G2430gat,G2431gat,G2432gat,G2435gat,G2436gat,G2437gat,G2438gat,G2439gat,G2440gat,G2443gat,G2444gat,G2445gat,G2448gat,G2449gat,G2450gat,G2467gat,G2468gat,G2469gat,G2470gat,G2471gat,G2474gat,G2475gat,G2476gat,G2477gat,G2478gat,G2481gat,G2482gat,G2483gat,G2486gat,G2487gat,G2632gat,G2633gat,G2634gat,G2635gat,G2636gat,G2637gat,G2638gat,G2639gat,G2640gat,G2641gat,G2642gat,G2643gat,G2644gat,G2645gat,G2646gat,G2647gat,G2648gat,G2652gat,G2656gat,G2659gat,G2662gat,G2666gat,G2670gat,G2673gat,G2677gat,G2681gat,G2684gat,G2688gat,G2692gat,G2697gat,G2702gat,G2706gat,G2710gat,G2715gat,G2719gat,G2723gat,G2728gat,G2729gat,G2730gat,G2731gat,G2732gat,G2733gat,G2734gat,G2735gat,G2736gat,G2737gat,G2738gat,G2739gat,G2740gat,G2741gat,G2742gat,G2743gat,G2744gat,G2745gat,G2746gat,G2748gat,G2749gat,G2750gat,G2751gat,G2754gat,G2755gat,G2756gat,G2757gat,G2758gat,G2761gat,G2764gat,G2768gat,G2769gat,G2898gat,G2899gat,G2900gat,G2901gat,G2962gat,G2966gat,G2967gat,G2973gat,G2977gat,G2980gat,G2984gat,G2985gat,G2986gat,G2987gat,G2988gat,G2989gat,G2990gat,G2991gat,G2992gat,G2993gat,G2994gat,G2995gat,G2996gat,G2997gat,G2998gat,G2999gat,G3000gat,G3001gat,G3002gat,G3003gat,G3004gat,G3005gat,G3006gat,G3007gat,G3008gat,G3009gat,G3010gat,G3011gat,G3012gat,G3013gat,G3014gat,G3015gat,G3016gat,G3017gat,G3018gat,G3019gat,G3020gat,G3021gat,G3022gat,G3023gat,G3024gat,G3025gat,G3026gat,G3027gat,G3028gat,G3029gat,G3030gat,G3031gat,G3032gat,G3033gat,G3034gat,G3035gat,G3036gat,G3037gat,G3038gat,G3039gat,G3040gat,G3041gat,G3042gat,G3043gat,G3044gat,G3045gat,G3046gat,G3047gat,G3048gat,G3049gat,G3050gat,G3051gat,G3052gat,G3053gat,G3054gat,G3055gat,G3056gat,G3057gat,G3058gat,G3059gat,G3060gat,G3061gat,G3062gat,G3063gat,G3064gat,G3065gat,G3066gat,G3067gat,G3068gat,G3069gat,G3070gat,G3071gat,G3072gat,G3073gat,G3074gat,G3075gat,G3076gat,G3077gat,G3078gat,G3079gat,G3080gat,G3081gat,G3082gat,G3083gat,G3084gat,G3085gat,G3086gat,G3087gat,G3088gat,G3089gat,G3090gat,G3091gat,G3092gat,G3093gat,G3094gat,G3095gat,G3096gat,G3097gat,G3098gat,G3099gat,G3100gat,G3101gat,G3102gat,G3103gat,G3104gat,G3105gat,G3106gat,G3107gat,G3108gat,G3109gat,G3110gat,G3111gat,G3115gat,G3118gat,G3119gat,G3125gat,G3131gat,G3134gat,G3138gat,G3141gat,G3145gat,G3148gat,G3149gat,G3155gat,G3161gat,G3164gat,G3168gat,G3171gat,G3172gat,G3175gat,G3178gat,G3181gat,G3184gat,G3187gat,G3190gat,G3191gat,G3192gat,G3193gat,G3194gat,G3196gat,G3206gat,G3207gat,G3208gat,G3209gat,G3210gat,G3211gat,G3212gat,G3213gat,G3214gat,G3215gat,G3216gat,G3217gat,G3218gat,G3219gat,G3220gat,G3221gat,G3222gat,G3223gat,G3224gat,G3225gat,G3226gat,G3227gat,G3228gat,G3229gat,G3230gat,G3231gat,G3232gat,G3233gat,G3234gat,G3235gat,G3236gat,G3237gat,G3238gat,G3239gat,G3240gat,G3241gat,G3242gat,G3243gat,G3244gat,G3245gat,G3246gat,G3247gat,G3248gat,G3249gat,G3250gat,G3251gat,G3252gat,G3253gat,G3254gat,G3255gat,G3256gat,G3257gat,G3258gat,G3259gat,G3260gat,G3261gat,G3262gat,G3263gat,G3264gat,G3265gat,G3266gat,G3267gat,G3268gat,G3269gat,G3270gat,G3271gat,G3272gat,G3273gat,G3274gat,G3275gat,G3276gat,G3277gat,G3278gat,G3279gat,G3280gat,G3281gat,G3282gat,G3283gat,G3284gat,G3285gat,G3286gat,G3287gat,G3288gat,G3289gat,G3290gat,G3291gat,G3292gat,G3293gat,G3294gat,G3295gat,G3296gat,G3297gat,G3298gat,G3299gat,G3300gat,G3301gat,G3302gat,G3303gat,G3304gat,G3305gat,G3306gat,G3307gat,G3308gat,G3309gat,G3310gat,G3311gat,G3312gat,G3313gat,G3314gat,G3315gat,G3316gat,G3317gat,G3318gat,G3319gat,G3320gat,G3321gat,G3322gat,G3323gat,G3324gat,G3325gat,G3326gat,G3327gat,G3328gat,G3329gat,G3330gat,G3331gat,G3332gat,G3333gat,G3334gat,G3383gat,G3387gat,G3388gat,G3389gat,G33890gat,G33891gat,G3390gat,G33900gat,G33901gat,G3391gat,G33910gat,G33911gat,G3392gat,G33920gat,G33921gat,G3393gat,G33930gat,G33931gat,G3394gat,G33940gat,G33941gat,G3395gat,G33950gat,G33951gat,G3396gat,G33960gat,G33961gat,G3397gat,G33970gat,G33971gat,G3398gat,G33980gat,G33981gat,G3399gat,G33990gat,G33991gat,G3400gat,G34000gat,G34001gat,G3401gat,G34010gat,G34011gat,G3402gat,G34020gat,G34021gat,G3403gat,G34030gat,G34031gat,G3404gat,G34040gat,G34041gat,G3405gat,G3406gat,G3407gat,G3410gat,G3413gat,G3414gat,G3415gat,G3419gat,G3423gat,G3426gat,G3429gat,G3430gat,G3431gat,G3434gat,G3437gat,G3438gat,G3439gat,G3442gat,G3445gat,G3446gat,G3447gat,G3451gat,G3455gat,G3458gat,G3461gat,G3462gat,G3463gat,G3466gat,G3469gat,G3470gat,G3471gat,G3534gat,G3535gat,G3536gat,G3537gat,G3538gat,G3539gat,G3540gat,G3541gat,G3542gat,G3543gat,G3544gat,G3545gat,G3546gat,G3547gat,G3548gat,G3549gat,G3550gat,G3551gat,G3552gat,G3557gat,G3568gat,G3573gat,G3578gat,G3589gat,G3594gat,G3605gat,G3626gat,G3627gat,G3628gat,G3629gat,G3630gat,G3631gat,G3632gat,G3633gat,G3634gat,G3635gat,G3636gat,G3637gat,G3638gat,G3639gat,G3640gat,G3641gat,G3642gat,G3643gat,G3644gat,G3645gat,G3648gat,G3651gat,G3652gat,G3653gat,G3654gat,G3657gat,G3658gat,G3661gat,G3662gat,G3663gat,G3664gat,G3667gat,G3670gat,G3671gat,G3672gat,G3673gat,G3676gat,G3677gat,G3680gat,G3681gat,G3682gat,G3685gat,G3686gat,G3687gat,G3688gat,G3689gat,G3690gat,G3693gat,G3694gat,G3695gat,G3696gat,G3703gat,G3704gat,G3705gat,G3706gat,G3707gat,G3708gat,G3711gat,G3712gat,G3713gat,G3714gat,G3715gat,G3716gat,G3717gat,G3718gat,G3719gat,G3720gat,G3721gat,G3731gat,G3734gat,G3740gat,G3743gat,G3753gat,G3756gat,G3762gat,G3765gat,G3766gat,G3773gat,G3774gat,G3775gat,G3776gat,G3777gat,G3778gat,G3779gat,G3780gat,G3786gat,G3789gat,G3800gat,G3803gat,G3809gat,G3812gat,G3815gat,G3818gat,G3834gat,G3835gat,G3838gat,G3845gat,G3884gat,G3885gat,G3894gat,G3895gat,G3898gat,G3899gat,G3906gat,G3911gat,G3912gat,G3916gat,G3920gat,G3924gat,G3925gat,G3926gat,G3930gat,G3931gat,G3932gat,G3935gat,G3936gat,G3947gat,G3948gat,G3992gat,G3996gat,G4013gat,G4029gat,G4030gat,G4031gat,G4032gat,G4033gat,G4034gat,G4042gat,G4043gat,G4044gat,G4045gat,G4046gat,G4047gat,G4048gat,G4049gat,G4050gat,G4051gat,G4052gat,G4053gat,G4054gat,G4055gat,G4056gat,G4057gat,G4058gat,G4065gat,G4066gat,G4073gat,G4074gat,G4075gat,G4076gat,G4077gat,G4078gat,G4079gat,G4080gat,G4085gat,G4086gat,G4088gat,G4090gat,G4091gat,G4094gat,G4098gat,G4101gat,G4104gat,G4105gat,G4106gat,G4107gat,G4108gat,G4109gat,G4110gat,G4111gat,G4112gat,G4113gat,G4114gat,G4115gat,G4116gat,G4119gat,G4122gat,G4123gat,G4126gat,G4127gat,G4128gat,G4139gat,G4142gat,G4146gat,G4147gat,G4148gat,G4149gat,G4150gat,G4151gat,G4152gat,G4153gat,G4154gat,G4161gat,G4186gat,G4189gat,G4190gat,G4191gat,G4192gat,G4193gat,G4194gat,G4195gat,G4196gat,G4197gat,G4218gat,G4238gat,G4239gat,G4241gat,G4242gat,G4251gat,G4252gat,G4253gat,G4254gat,G4255gat,G4256gat,G4257gat,G4258gat,G4283gat,G4284gat,G4287gat,G4291gat,G4295gat,G4299gat,G4303gat,G4304gat,G4310gat,G4316gat,G4317gat,G4318gat,G4319gat,G4322gat,G4325gat,G4326gat,G4327gat,G4328gat,G4329gat,G4330gat,G4331gat,G4335gat,G4338gat,G4341gat,G4344gat,G4347gat,G4350gat,G4371gat,G4376gat,G4377gat,G4387gat,G4390gat,G4393gat,G4416gat,G4421gat,G4427gat,G4435gat,G4442gat,G4443gat,G4446gat,G4447gat,G4448gat,G4452gat,G4458gat,G4461gat,G4462gat,G4463gat,G4464gat,G4468gat,G4472gat,G4475gat,G4484gat,G4486gat,G4487gat,G4491gat,G4493gat,G4496gat,G4497gat,G4498gat,G4503gat,G4506gat,G4507gat,G4508gat,G4509gat,G4510gat,G4511gat,G4515gat,G4526gat,G4527gat,G4528gat,G4529gat,G4530gat,G4545gat,G4549gat,G4552gat,G4555gat,G4558gat,G4559gat,G4562gat,G4563gat,G4568gat,G4572gat,G4573gat,G4576gat,G4587gat,G4588gat,G4593gat,G4596gat,G4597gat,G4599gat,G4602gat,G4603gat,G4608gat,G4619gat,G4623gat,G4628gat,G4629gat,G4630gat,G4635gat,G4636gat,G4640gat,G4641gat,G4642gat,G4643gat,G4644gat,G4647gat,G4650gat,G4668gat,G4669gat,G4670gat,G4673gat,G4674gat,G4675gat,G4676gat,G4677gat,G4678gat,G4679gat,G4687gat,G4688gat,G4704gat,G4705gat,G4706gat,G4707gat,G4708gat,G4711gat,G4716gat,G4717gat,G4721gat,G4726gat,G4727gat,G4730gat,G4733gat,G4740gat,G4743gat,G4747gat,G4748gat,G4749gat,G4750gat,G4753gat,G4754gat,G4755gat,G4756gat,G4757gat,G4769gat,G4772gat,G4775gat,G4778gat,G4786gat,G4787gat,G4788gat,G4789gat,G4794gat,G4797gat,G4800gat,G4808gat,G4816gat,G4817gat,G4818gat,G4822gat,G4823gat,G4826gat,G4829gat,G4830gat,G4831gat,G4838gat,G4859gat,G4860gat,G4868gat,G4870gat,G4872gat,G4873gat,G4876gat,G4880gat,G4885gat,G4889gat,G4895gat,G4896gat,G4897gat,G4898gat,G4899gat,G4900gat,G4901gat,G4902gat,G4904gat,G4905gat,G4906gat,G4907gat,G4913gat,G4916gat,G4920gat,G4921gat,G4924gat,G4925gat,G4926gat,G4928gat,G4929gat,G4930gat,G4931gat,G4946gat,G4949gat,G4950gat,G4951gat,G4952gat,G4953gat,G4954gat,G4957gat,G4964gat,G4965gat,G4968gat,G4969gat,G4970gat,G4973gat,G4978gat,G4979gat,G4980gat,G4981gat,G4982gat,G4983gat,G4984gat,G4985gat,G4988gat,G4991gat,G4996gat,G4999gat,G5007gat,G5010gat,G5013gat,G5018gat,G5021gat,G5026gat,G5029gat,G5030gat,G5046gat,G5050gat,G5055gat,G5058gat,G5061gat,G5066gat,G5080gat,G5085gat,G5094gat,G5095gat,G5097gat,G5103gat,G5108gat,G5109gat,G5110gat,G5114gat,G5122gat,G5125gat,G5128gat,G5133gat,G5136gat,G5145gat,G5159gat,G5166gat,G5173gat,G5182gat,G5183gat,G5193gat,G5196gat,G5197gat,G5198gat,G5199gat,G5201gat,G5203gat,G5212gat,G5215gat,G5217gat,G5219gat,G5220gat,G5221gat,G5222gat,G5223gat,G5224gat,G5225gat,G5228gat,G5232gat,G5233gat,G5234gat,G5235gat,G5236gat,G5240gat,G5242gat,G5243gat,G5245gat,G5246gat,G5250gat,G5253gat,G5254gat,G5257gat,G5258gat,G5261gat,G5266gat,G5277gat,G5278gat,G5279gat,G5283gat,G5284gat,G5285gat,G5286gat,G5295gat,G5298gat,G5309gat,G5312gat,G5313gat,G5322gat,G5323gat,G5340gat,G5341gat,G5344gat,G5345gat,G5348gat,G5349gat,G5350gat,G5351gat,G5352gat,G5353gat,G5354gat,G5355gat,G5356gat,G5357gat,G5358gat,G5359gat,G5361gat_enc,nXOR0,nXOR1,nXOR2,nXOR3,nXOR4,nXOR5,nXOR6,nXOR7,not_keyinp0,not_keyinp1,not_keyinp2,not_keyinp3,not_keyinp4,not_keyinp5,not_keyinp6,not_keyinp7,flipSig,maskSig,not_mask,flip_mask;

not NOT1_1 (G665gat, G50gat);
not NOT1_2 (G679gat, G58gat);
not NOT1_3 (G686gat, G68gat);
not NOT1_4 (G702gat, G77gat);
not NOT1_5 (G724gat, G87gat);
not NOT1_6 (G736gat, G97gat);
not NOT1_7 (G749gat, G107gat);
not NOT1_8 (G763gat, G116gat);
or OR2_9 (G768gat, G257gat, G264gat);
not NOT1_10 (G769gat, G1gat);
not NOT1_11 (G779gat, G1gat);
not NOT1_12 (G786gat, G13gat);
and AND2_13 (G793gat, G13gat, G20gat);
not NOT1_14 (G794gat, G20gat);
not NOT1_15 (G803gat, G20gat);
not NOT1_16 (G820gat, G33gat);
not NOT1_17 (G825gat, G33gat);
and AND2_18 (G829gat, G33gat, G41gat);
not NOT1_19 (G832gat, G41gat);
or OR2_20 (G835gat, G41gat, G45gat);
not NOT1_21 (G839gat, G45gat);
not NOT1_22 (G842gat, G50gat);
not NOT1_23 (G848gat, G58gat);
not NOT1_24 (G854gat, G68gat);
not NOT1_25 (G861gat, G87gat);
not NOT1_26 (G867gat, G97gat);
not NOT1_27 (G870gat, G107gat);
not NOT1_28 (G883gat, G20gat);
not NOT1_29 (G889gat, G200gat);
and AND2_30 (G890gat, G20gat, G200gat);
nand NAND2_31 (G891gat, G20gat, G200gat);
and AND2_32 (G892gat, G20gat, G179gat);
not NOT1_33 (G895gat, G20gat);
or OR2_34 (G896gat, G349gat, G33gat);
nand NAND2_35 (G913gat, G1gat, G13gat);
nand NAND3_36 (G914gat, G1gat, G20gat, G33gat);
not NOT1_37 (G915gat, G20gat);
not NOT1_38 (G916gat, G33gat);
not NOT1_39 (G920gat, G213gat);
and AND2_40 (G1067gat, G250gat, G768gat);
or OR2_41 (G1117gat, G820gat, G20gat);
or OR2_42 (G1179gat, G895gat, G169gat);
not NOT1_43 (G1196gat, G793gat);
or OR2_44 (G1197gat, G915gat, G1gat);
and AND2_45 (G1202gat, G913gat, G914gat);
or OR2_46 (G1219gat, G916gat, G1gat);
and AND3_47 (G1250gat, G842gat, G848gat, G854gat);
nand NAND2_48 (G1251gat, G226gat, G655gat);
nand NAND2_49 (G1252gat, G232gat, G670gat);
nand NAND2_50 (G1253gat, G238gat, G690gat);
nand NAND2_51 (G1254gat, G244gat, G706gat);
nand NAND2_52 (G1255gat, G250gat, G715gat);
nand NAND2_53 (G1256gat, G257gat, G727gat);
nand NAND2_54 (G1257gat, G264gat, G740gat);
nand NAND2_55 (G1258gat, G270gat, G753gat);
not NOT1_56 (G1259gat, G926gat);
not NOT1_57 (G1260gat, G929gat);
not NOT1_58 (G1261gat, G932gat);
not NOT1_59 (G1262gat, G935gat);
nand NAND2_60 (G1263gat, G679gat, G686gat);
nand NAND2_61 (G1264gat, G736gat, G749gat);
nand NAND2_62 (G1267gat, G683gat, G699gat);
not NOT1_63 (G1271gat, G953gat);
not NOT1_64 (G1272gat, G959gat);
and AND2_65 (G1306gat, G779gat, G835gat);
and AND3_66 (G1315gat, G779gat, G836gat, G832gat);
and AND2_67 (G1322gat, G769gat, G836gat);
and AND3_68 (G1325gat, G772gat, G786gat, G798gat);
nand NAND3_69 (G1328gat, G772gat, G786gat, G798gat);
nand NAND2_70 (G1331gat, G772gat, G786gat);
nand NAND3_71 (G1337gat, G782gat, G794gat, G45gat);
nand NAND3_72 (G1338gat, G842gat, G848gat, G854gat);
not NOT1_73 (G1339gat, G956gat);
and AND3_74 (G1340gat, G861gat, G867gat, G870gat);
nand NAND3_75 (G1343gat, G861gat, G867gat, G870gat);
not NOT1_76 (G1344gat, G962gat);
not NOT1_77 (G1345gat, G803gat);
not NOT1_78 (G1346gat, G803gat);
not NOT1_79 (G1347gat, G803gat);
not NOT1_80 (G1348gat, G803gat);
not NOT1_81 (G1349gat, G803gat);
not NOT1_82 (G1350gat, G803gat);
not NOT1_83 (G1351gat, G803gat);
not NOT1_84 (G1352gat, G803gat);
or OR2_85 (G1353gat, G883gat, G886gat);
nor NOR2_86 (G1358gat, G883gat, G886gat);
not NOT1_87 (G1366gat, G892gat);
not NOT1_88 (G1401gat, G896gat);
not NOT1_89 (G1402gat, G896gat);
not NOT1_90 (G1403gat, G896gat);
not NOT1_91 (G1404gat, G896gat);
not NOT1_92 (G1405gat, G896gat);
not NOT1_93 (G1406gat, G896gat);
not NOT1_94 (G1407gat, G896gat);
not NOT1_95 (G1408gat, G896gat);
or OR2_96 (G1409gat, G1gat, G1196gat);
not NOT1_97 (G1426gat, G829gat);
not NOT1_98 (G1427gat, G829gat);
and AND3_99 (G1452gat, G769gat, G782gat, G794gat);
not NOT1_100 (G1459gat, G917gat);
not NOT1_101 (G1460gat, G965gat);
or OR2_102 (G1461gat, G920gat, G923gat);
nor NOR2_103 (G1464gat, G920gat, G923gat);
not NOT1_104 (G1467gat, G938gat);
not NOT1_105 (G1468gat, G941gat);
not NOT1_106 (G1469gat, G944gat);
not NOT1_107 (G1470gat, G947gat);
not NOT1_108 (G1474gat, G950gat);
nand NAND2_109 (G1505gat, G702gat, G1250gat);
and AND4_110 (G1507gat, G1251gat, G1252gat, G1253gat, G1254gat);
and AND4_111 (G1508gat, G1255gat, G1256gat, G1257gat, G1258gat);
nand NAND2_112 (G1509gat, G929gat, G1259gat);
nand NAND2_113 (G1510gat, G926gat, G1260gat);
nand NAND2_114 (G1511gat, G935gat, G1261gat);
nand NAND2_115 (G1512gat, G932gat, G1262gat);
and AND2_116 (G1520gat, G655gat, G1263gat);
and AND2_117 (G1562gat, G874gat, G1337gat);
not NOT1_118 (G1579gat, G1117gat);
and AND2_119 (G1580gat, G803gat, G1117gat);
and AND2_120 (G1581gat, G1338gat, G1345gat);
not NOT1_121 (G1582gat, G1117gat);
and AND2_122 (G1583gat, G803gat, G1117gat);
not NOT1_123 (G1584gat, G1117gat);
and AND2_124 (G1585gat, G803gat, G1117gat);
and AND2_125 (G1586gat, G854gat, G1347gat);
not NOT1_126 (G1587gat, G1117gat);
and AND2_127 (G1588gat, G803gat, G1117gat);
and AND2_128 (G1589gat, G77gat, G1348gat);
not NOT1_129 (G1590gat, G1117gat);
and AND2_130 (G1591gat, G803gat, G1117gat);
and AND2_131 (G1592gat, G1343gat, G1349gat);
not NOT1_132 (G1593gat, G1117gat);
and AND2_133 (G1594gat, G803gat, G1117gat);
not NOT1_134 (G1595gat, G1117gat);
and AND2_135 (G1596gat, G803gat, G1117gat);
and AND2_136 (G1597gat, G870gat, G1351gat);
not NOT1_137 (G1598gat, G1117gat);
and AND2_138 (G1599gat, G803gat, G1117gat);
and AND2_139 (G1600gat, G116gat, G1352gat);
and AND2_140 (G1643gat, G222gat, G1401gat);
and AND2_141 (G1644gat, G223gat, G1402gat);
and AND2_142 (G1645gat, G226gat, G1403gat);
and AND2_143 (G1646gat, G232gat, G1404gat);
and AND2_144 (G1647gat, G238gat, G1405gat);
and AND2_145 (G1648gat, G244gat, G1406gat);
and AND2_146 (G1649gat, G250gat, G1407gat);
and AND2_147 (G1650gat, G257gat, G1408gat);
and AND3_148 (G1667gat, G1gat, G13gat, G1426gat);
and AND3_149 (G1670gat, G1gat, G13gat, G1427gat);
not NOT1_150 (G1673gat, G1202gat);
not NOT1_151 (G1674gat, G1202gat);
not NOT1_152 (G1675gat, G1202gat);
not NOT1_153 (G1676gat, G1202gat);
not NOT1_154 (G1677gat, G1202gat);
not NOT1_155 (G1678gat, G1202gat);
not NOT1_156 (G1679gat, G1202gat);
not NOT1_157 (G1680gat, G1202gat);
nand NAND2_158 (G1691gat, G941gat, G1467gat);
nand NAND2_159 (G1692gat, G938gat, G1468gat);
nand NAND2_160 (G1693gat, G947gat, G1469gat);
nand NAND2_161 (G1694gat, G944gat, G1470gat);
not NOT1_162 (G1713gat, G1505gat);
and AND2_163 (G1714gat, G87gat, G1264gat);
nand NAND2_164 (G1715gat, G1509gat, G1510gat);
nand NAND2_165 (G1718gat, G1511gat, G1512gat);
nand NAND2_166 (G1721gat, G1507gat, G1508gat);
and AND2_167 (G1722gat, G763gat, G1340gat);
nand NAND2_168 (G1725gat, G763gat, G1340gat);
not NOT1_169 (G1726gat, G1268gat);
nand NAND2_170 (G1727gat, G1493gat, G1271gat);
not NOT1_171 (G1728gat, G1493gat);
and AND2_172 (G1729gat, G683gat, G1268gat);
nand NAND2_173 (G1730gat, G1499gat, G1272gat);
not NOT1_174 (G1731gat, G1499gat);
nand NAND2_175 (G1735gat, G87gat, G1264gat);
not NOT1_176 (G1736gat, G1273gat);
not NOT1_177 (G1737gat, G1276gat);
nand NAND2_178 (G1738gat, G1325gat, G821gat);
nand NAND2_179 (G1747gat, G1325gat, G825gat);
nand NAND3_180 (G1756gat, G772gat, G1279gat, G798gat);
nand NAND4_181 (G1761gat, G772gat, G786gat, G798gat, G1302gat);
nand NAND2_182 (G1764gat, G1496gat, G1339gat);
not NOT1_183 (G1765gat, G1496gat);
nand NAND2_184 (G1766gat, G1502gat, G1344gat);
not NOT1_185 (G1767gat, G1502gat);
not NOT1_186 (G1768gat, G1328gat);
not NOT1_187 (G1769gat, G1334gat);
not NOT1_188 (G1770gat, G1331gat);
and AND2_189 (G1787gat, G845gat, G1579gat);
and AND2_190 (G1788gat, G150gat, G1580gat);
and AND2_191 (G1789gat, G851gat, G1582gat);
and AND2_192 (G1790gat, G159gat, G1583gat);
and AND2_193 (G1791gat, G77gat, G1584gat);
and AND2_194 (G1792gat, G50gat, G1585gat);
and AND2_195 (G1793gat, G858gat, G1587gat);
and AND2_196 (G1794gat, G845gat, G1588gat);
and AND2_197 (G1795gat, G864gat, G1590gat);
and AND2_198 (G1796gat, G851gat, G1591gat);
and AND2_199 (G1797gat, G107gat, G1593gat);
and AND2_200 (G1798gat, G77gat, G1594gat);
and AND2_201 (G1799gat, G116gat, G1595gat);
and AND2_202 (G1800gat, G858gat, G1596gat);
and AND2_203 (G1801gat, G283gat, G1598gat);
and AND2_204 (G1802gat, G864gat, G1599gat);
and AND2_205 (G1803gat, G200gat, G1363gat);
and AND2_206 (G1806gat, G889gat, G1363gat);
and AND2_207 (G1809gat, G890gat, G1366gat);
and AND2_208 (G1812gat, G891gat, G1366gat);
nand NAND2_209 (G1815gat, G1298gat, G1302gat);
nand NAND2_210 (G1818gat, G821gat, G1302gat);
nand NAND3_211 (G1821gat, G772gat, G1279gat, G1179gat);
nand NAND3_212 (G1824gat, G786gat, G794gat, G1298gat);
nand NAND2_213 (G1833gat, G786gat, G1298gat);
not NOT1_214 (G1842gat, G1369gat);
not NOT1_215 (G1843gat, G1369gat);
not NOT1_216 (G1844gat, G1369gat);
not NOT1_217 (G1845gat, G1369gat);
not NOT1_218 (G1846gat, G1369gat);
not NOT1_219 (G1847gat, G1369gat);
not NOT1_220 (G1848gat, G1369gat);
not NOT1_221 (G1849gat, G1384gat);
and AND2_222 (G1850gat, G1384gat, G896gat);
not NOT1_223 (G1851gat, G1384gat);
and AND2_224 (G1852gat, G1384gat, G896gat);
not NOT1_225 (G1853gat, G1384gat);
and AND2_226 (G1854gat, G1384gat, G896gat);
not NOT1_227 (G1855gat, G1384gat);
and AND2_228 (G1856gat, G1384gat, G896gat);
not NOT1_229 (G1857gat, G1384gat);
and AND2_230 (G1858gat, G1384gat, G896gat);
not NOT1_231 (G1859gat, G1384gat);
and AND2_232 (G1860gat, G1384gat, G896gat);
not NOT1_233 (G1861gat, G1384gat);
and AND2_234 (G1862gat, G1384gat, G896gat);
not NOT1_235 (G1863gat, G1384gat);
and AND2_236 (G1864gat, G1384gat, G896gat);
and AND2_237 (G1869gat, G1202gat, G1409gat);
nor NOR2_238 (G1870gat, G50gat, G1409gat);
not NOT1_239 (G1873gat, G1306gat);
and AND2_240 (G1874gat, G1202gat, G1409gat);
nor NOR2_241 (G1875gat, G58gat, G1409gat);
not NOT1_242 (G1878gat, G1306gat);
and AND2_243 (G1879gat, G1202gat, G1409gat);
nor NOR2_244 (G1880gat, G68gat, G1409gat);
not NOT1_245 (G1883gat, G1306gat);
and AND2_246 (G1884gat, G1202gat, G1409gat);
nor NOR2_247 (G1885gat, G77gat, G1409gat);
not NOT1_248 (G1888gat, G1306gat);
and AND2_249 (G1889gat, G1202gat, G1409gat);
nor NOR2_250 (G1890gat, G87gat, G1409gat);
not NOT1_251 (G1893gat, G1322gat);
and AND2_252 (G1894gat, G1202gat, G1409gat);
nor NOR2_253 (G1895gat, G97gat, G1409gat);
not NOT1_254 (G1898gat, G1315gat);
and AND2_255 (G1899gat, G1202gat, G1409gat);
nor NOR2_256 (G1900gat, G107gat, G1409gat);
not NOT1_257 (G1903gat, G1315gat);
and AND2_258 (G1904gat, G1202gat, G1409gat);
nor NOR2_259 (G1905gat, G116gat, G1409gat);
not NOT1_260 (G1908gat, G1315gat);
and AND2_261 (G1909gat, G1452gat, G213gat);
nand NAND2_262 (G1912gat, G1452gat, G213gat);
and AND3_263 (G1913gat, G1452gat, G213gat, G343gat);
nand NAND3_264 (G1917gat, G1452gat, G213gat, G343gat);
and AND3_265 (G1922gat, G1452gat, G213gat, G343gat);
nand NAND3_266 (G1926gat, G1452gat, G213gat, G343gat);
nand NAND2_267 (G1933gat, G1691gat, G1692gat);
nand NAND2_268 (G1936gat, G1693gat, G1694gat);
not NOT1_269 (G1939gat, G1471gat);
nand NAND2_270 (G1940gat, G1471gat, G1474gat);
not NOT1_271 (G1941gat, G1475gat);
not NOT1_272 (G1942gat, G1478gat);
not NOT1_273 (G1943gat, G1481gat);
not NOT1_274 (G1944gat, G1484gat);
not NOT1_275 (G1945gat, G1487gat);
not NOT1_276 (G1946gat, G1490gat);
not NOT1_277 (G1947gat, G1714gat);
nand NAND2_278 (G1960gat, G953gat, G1728gat);
nand NAND2_279 (G1961gat, G959gat, G1731gat);
and AND2_280 (G1966gat, G1520gat, G1276gat);
nand NAND2_281 (G1981gat, G956gat, G1765gat);
nand NAND2_282 (G1982gat, G962gat, G1767gat);
and AND2_283 (G1983gat, G1067gat, G1768gat);
or OR3_284 (G1986gat, G1581gat, G1787gat, G1788gat);
or OR3_285 (G1987gat, G1586gat, G1791gat, G1792gat);
or OR3_286 (G1988gat, G1589gat, G1793gat, G1794gat);
or OR3_287 (G1989gat, G1592gat, G1795gat, G1796gat);
or OR3_288 (G1990gat, G1597gat, G1799gat, G1800gat);
or OR3_289 (G1991gat, G1600gat, G1801gat, G1802gat);
and AND2_290 (G2022gat, G77gat, G1849gat);
and AND2_291 (G2023gat, G223gat, G1850gat);
and AND2_292 (G2024gat, G87gat, G1851gat);
and AND2_293 (G2025gat, G226gat, G1852gat);
and AND2_294 (G2026gat, G97gat, G1853gat);
and AND2_295 (G2027gat, G232gat, G1854gat);
and AND2_296 (G2028gat, G107gat, G1855gat);
and AND2_297 (G2029gat, G238gat, G1856gat);
and AND2_298 (G2030gat, G116gat, G1857gat);
and AND2_299 (G2031gat, G244gat, G1858gat);
and AND2_300 (G2032gat, G283gat, G1859gat);
and AND2_301 (G2033gat, G250gat, G1860gat);
and AND2_302 (G2034gat, G294gat, G1861gat);
and AND2_303 (G2035gat, G257gat, G1862gat);
and AND2_304 (G2036gat, G303gat, G1863gat);
and AND2_305 (G2037gat, G264gat, G1864gat);
not NOT1_306 (G2043gat, G1667gat);
not NOT1_307 (G2057gat, G1670gat);
and AND3_308 (G2068gat, G50gat, G1197gat, G1869gat);
and AND3_309 (G2073gat, G58gat, G1197gat, G1874gat);
and AND3_310 (G2078gat, G68gat, G1197gat, G1879gat);
and AND3_311 (G2083gat, G77gat, G1197gat, G1884gat);
and AND3_312 (G2088gat, G87gat, G1219gat, G1889gat);
and AND3_313 (G2093gat, G97gat, G1219gat, G1894gat);
and AND3_314 (G2098gat, G107gat, G1219gat, G1899gat);
and AND3_315 (G2103gat, G116gat, G1219gat, G1904gat);
not NOT1_316 (G2121gat, G1562gat);
not NOT1_317 (G2122gat, G1562gat);
not NOT1_318 (G2123gat, G1562gat);
not NOT1_319 (G2124gat, G1562gat);
not NOT1_320 (G2125gat, G1562gat);
not NOT1_321 (G2126gat, G1562gat);
not NOT1_322 (G2127gat, G1562gat);
not NOT1_323 (G2128gat, G1562gat);
nand NAND2_324 (G2133gat, G950gat, G1939gat);
nand NAND2_325 (G2134gat, G1478gat, G1941gat);
nand NAND2_326 (G2135gat, G1475gat, G1942gat);
nand NAND2_327 (G2136gat, G1484gat, G1943gat);
nand NAND2_328 (G2137gat, G1481gat, G1944gat);
nand NAND2_329 (G2138gat, G1490gat, G1945gat);
nand NAND2_330 (G2139gat, G1487gat, G1946gat);
not NOT1_331 (G2141gat, G1933gat);
not NOT1_332 (G2142gat, G1936gat);
not NOT1_333 (G2143gat, G1738gat);
and AND2_334 (G2144gat, G1738gat, G1747gat);
not NOT1_335 (G2145gat, G1747gat);
nand NAND2_336 (G2146gat, G1727gat, G1960gat);
nand NAND2_337 (G2147gat, G1730gat, G1961gat);
and AND4_338 (G2148gat, G1722gat, G1267gat, G665gat, G58gat);
not NOT1_339 (G2149gat, G1738gat);
and AND2_340 (G2150gat, G1738gat, G1747gat);
not NOT1_341 (G2151gat, G1747gat);
not NOT1_342 (G2152gat, G1738gat);
not NOT1_343 (G2153gat, G1747gat);
and AND2_344 (G2154gat, G1738gat, G1747gat);
not NOT1_345 (G2155gat, G1738gat);
not NOT1_346 (G2156gat, G1747gat);
and AND2_347 (G2157gat, G1738gat, G1747gat);
nand NAND2_348 (G2178gat, G1764gat, G1981gat);
nand NAND2_349 (G2179gat, G1766gat, G1982gat);
not NOT1_350 (G2180gat, G1756gat);
and AND2_351 (G2181gat, G1756gat, G1328gat);
not NOT1_352 (G2183gat, G1756gat);
and AND2_353 (G2184gat, G1331gat, G1756gat);
nand NAND2_354 (G2185gat, G1358gat, G1812gat);
nand NAND2_355 (G2188gat, G1358gat, G1809gat);
nand NAND2_356 (G2191gat, G1353gat, G1812gat);
nand NAND2_357 (G2194gat, G1353gat, G1809gat);
nand NAND2_358 (G2197gat, G1358gat, G1806gat);
nand NAND2_359 (G2200gat, G1358gat, G1803gat);
nand NAND2_360 (G2203gat, G1353gat, G1806gat);
nand NAND2_361 (G2206gat, G1353gat, G1803gat);
not NOT1_362 (G2209gat, G1815gat);
not NOT1_363 (G2210gat, G1818gat);
and AND2_364 (G2211gat, G1815gat, G1818gat);
not NOT1_365 (G2230gat, G1833gat);
not NOT1_366 (G2231gat, G1833gat);
not NOT1_367 (G2232gat, G1833gat);
not NOT1_368 (G2233gat, G1833gat);
not NOT1_369 (G2234gat, G1824gat);
not NOT1_370 (G2235gat, G1824gat);
not NOT1_371 (G2236gat, G1824gat);
not NOT1_372 (G2237gat, G1824gat);
or OR3_373 (G2238gat, G2022gat, G1643gat, G2023gat);
or OR3_374 (G2239gat, G2024gat, G1644gat, G2025gat);
or OR3_375 (G2240gat, G2026gat, G1645gat, G2027gat);
or OR3_376 (G2241gat, G2028gat, G1646gat, G2029gat);
or OR3_377 (G2242gat, G2030gat, G1647gat, G2031gat);
or OR3_378 (G2243gat, G2032gat, G1648gat, G2033gat);
or OR3_379 (G2244gat, G2034gat, G1649gat, G2035gat);
or OR3_380 (G2245gat, G2036gat, G1650gat, G2037gat);
and AND2_381 (G2270gat, G1986gat, G1673gat);
and AND2_382 (G2277gat, G1987gat, G1675gat);
and AND2_383 (G2282gat, G1988gat, G1676gat);
and AND2_384 (G2287gat, G1989gat, G1677gat);
and AND2_385 (G2294gat, G1990gat, G1679gat);
and AND2_386 (G2299gat, G1991gat, G1680gat);
and AND2_387 (G2307gat, G1930gat, G350gat);
nand NAND2_388 (G2310gat, G1930gat, G350gat);
nand NAND2_389 (G2325gat, G1940gat, G2133gat);
nand NAND2_390 (G2328gat, G2134gat, G2135gat);
nand NAND2_391 (G2331gat, G2136gat, G2137gat);
nand NAND2_392 (G2334gat, G2138gat, G2139gat);
nand NAND2_393 (G2341gat, G1936gat, G2141gat);
nand NAND2_394 (G2342gat, G1933gat, G2142gat);
and AND2_395 (G2347gat, G724gat, G2144gat);
and AND3_396 (G2348gat, G2146gat, G699gat, G1726gat);
and AND2_397 (G2349gat, G753gat, G2147gat);
and AND2_398 (G2350gat, G2148gat, G1273gat);
and AND2_399 (G2351gat, G736gat, G2150gat);
and AND2_400 (G2352gat, G1735gat, G2153gat);
and AND2_401 (G2353gat, G763gat, G2154gat);
and AND2_402 (G2354gat, G1725gat, G2156gat);
and AND2_403 (G2355gat, G749gat, G2157gat);
not NOT1_404 (G2374gat, G2178gat);
not NOT1_405 (G2375gat, G2179gat);
and AND2_406 (G2376gat, G1520gat, G2180gat);
and AND2_407 (G2379gat, G1721gat, G2181gat);
and AND2_408 (G2398gat, G665gat, G2211gat);
and AND3_409 (G2417gat, G2057gat, G226gat, G1873gat);
and AND3_410 (G2418gat, G2057gat, G274gat, G1306gat);
and AND2_411 (G2419gat, G2052gat, G2238gat);
and AND3_412 (G2420gat, G2057gat, G232gat, G1878gat);
and AND3_413 (G2421gat, G2057gat, G274gat, G1306gat);
and AND2_414 (G2422gat, G2052gat, G2239gat);
and AND3_415 (G2425gat, G2057gat, G238gat, G1883gat);
and AND3_416 (G2426gat, G2057gat, G274gat, G1306gat);
and AND2_417 (G2427gat, G2052gat, G2240gat);
and AND3_418 (G2430gat, G2057gat, G244gat, G1888gat);
and AND3_419 (G2431gat, G2057gat, G274gat, G1306gat);
and AND2_420 (G2432gat, G2052gat, G2241gat);
and AND3_421 (G2435gat, G2043gat, G250gat, G1893gat);
and AND3_422 (G2436gat, G2043gat, G274gat, G1322gat);
and AND2_423 (G2437gat, G2038gat, G2242gat);
and AND3_424 (G2438gat, G2043gat, G257gat, G1898gat);
and AND3_425 (G2439gat, G2043gat, G274gat, G1315gat);
and AND2_426 (G2440gat, G2038gat, G2243gat);
and AND3_427 (G2443gat, G2043gat, G264gat, G1903gat);
and AND3_428 (G2444gat, G2043gat, G274gat, G1315gat);
and AND2_429 (G2445gat, G2038gat, G2244gat);
and AND3_430 (G2448gat, G2043gat, G270gat, G1908gat);
and AND3_431 (G2449gat, G2043gat, G274gat, G1315gat);
and AND2_432 (G2450gat, G2038gat, G2245gat);
not NOT1_433 (G2467gat, G2313gat);
not NOT1_434 (G2468gat, G2316gat);
not NOT1_435 (G2469gat, G2319gat);
not NOT1_436 (G2470gat, G2322gat);
nand NAND2_437 (G2471gat, G2341gat, G2342gat);
not NOT1_438 (G2474gat, G2325gat);
not NOT1_439 (G2475gat, G2328gat);
not NOT1_440 (G2476gat, G2331gat);
not NOT1_441 (G2477gat, G2334gat);
or OR2_442 (G2478gat, G2348gat, G1729gat);
not NOT1_443 (G2481gat, G2175gat);
and AND2_444 (G2482gat, G2175gat, G1334gat);
and AND2_445 (G2483gat, G2349gat, G2183gat);
and AND2_446 (G2486gat, G2374gat, G1346gat);
and AND2_447 (G2487gat, G2375gat, G1350gat);
not NOT1_448 (G2632gat, G2212gat);
and AND2_449 (G2633gat, G2212gat, G1833gat);
not NOT1_450 (G2634gat, G2212gat);
and AND2_451 (G2635gat, G2212gat, G1833gat);
not NOT1_452 (G2636gat, G2212gat);
and AND2_453 (G2637gat, G2212gat, G1833gat);
not NOT1_454 (G2638gat, G2212gat);
and AND2_455 (G2639gat, G2212gat, G1833gat);
not NOT1_456 (G2640gat, G2221gat);
and AND2_457 (G2641gat, G2221gat, G1824gat);
not NOT1_458 (G2642gat, G2221gat);
and AND2_459 (G2643gat, G2221gat, G1824gat);
not NOT1_460 (G2644gat, G2221gat);
and AND2_461 (G2645gat, G2221gat, G1824gat);
not NOT1_462 (G2646gat, G2221gat);
and AND2_463 (G2647gat, G2221gat, G1824gat);
or OR3_464 (G2648gat, G2270gat, G1870gat, G2068gat);
nor NOR3_465 (G2652gat, G2270gat, G1870gat, G2068gat);
or OR3_466 (G2656gat, G2417gat, G2418gat, G2419gat);
or OR3_467 (G2659gat, G2420gat, G2421gat, G2422gat);
or OR3_468 (G2662gat, G2277gat, G1880gat, G2078gat);
nor NOR3_469 (G2666gat, G2277gat, G1880gat, G2078gat);
or OR3_470 (G2670gat, G2425gat, G2426gat, G2427gat);
or OR3_471 (G2673gat, G2282gat, G1885gat, G2083gat);
nor NOR3_472 (G2677gat, G2282gat, G1885gat, G2083gat);
or OR3_473 (G2681gat, G2430gat, G2431gat, G2432gat);
or OR3_474 (G2684gat, G2287gat, G1890gat, G2088gat);
nor NOR3_475 (G2688gat, G2287gat, G1890gat, G2088gat);
or OR3_476 (G2692gat, G2435gat, G2436gat, G2437gat);
or OR3_477 (G2697gat, G2438gat, G2439gat, G2440gat);
or OR3_478 (G2702gat, G2294gat, G1900gat, G2098gat);
nor NOR3_479 (G2706gat, G2294gat, G1900gat, G2098gat);
or OR3_480 (G2710gat, G2443gat, G2444gat, G2445gat);
or OR3_481 (G2715gat, G2299gat, G1905gat, G2103gat);
nor NOR3_482 (G2719gat, G2299gat, G1905gat, G2103gat);
or OR3_483 (G2723gat, G2448gat, G2449gat, G2450gat);
not NOT1_484 (G2728gat, G2304gat);
not NOT1_485 (G2729gat, G2158gat);
and AND2_486 (G2730gat, G1562gat, G2158gat);
not NOT1_487 (G2731gat, G2158gat);
and AND2_488 (G2732gat, G1562gat, G2158gat);
not NOT1_489 (G2733gat, G2158gat);
and AND2_490 (G2734gat, G1562gat, G2158gat);
not NOT1_491 (G2735gat, G2158gat);
and AND2_492 (G2736gat, G1562gat, G2158gat);
not NOT1_493 (G2737gat, G2158gat);
and AND2_494 (G2738gat, G1562gat, G2158gat);
not NOT1_495 (G2739gat, G2158gat);
and AND2_496 (G2740gat, G1562gat, G2158gat);
not NOT1_497 (G2741gat, G2158gat);
and AND2_498 (G2742gat, G1562gat, G2158gat);
not NOT1_499 (G2743gat, G2158gat);
and AND2_500 (G2744gat, G1562gat, G2158gat);
or OR3_501 (G2745gat, G2376gat, G1983gat, G2379gat);
nor NOR3_502 (G2746gat, G2376gat, G1983gat, G2379gat);
nand NAND2_503 (G2748gat, G2316gat, G2467gat);
nand NAND2_504 (G2749gat, G2313gat, G2468gat);
nand NAND2_505 (G2750gat, G2322gat, G2469gat);
nand NAND2_506 (G2751gat, G2319gat, G2470gat);
nand NAND2_507 (G2754gat, G2328gat, G2474gat);
nand NAND2_508 (G2755gat, G2325gat, G2475gat);
nand NAND2_509 (G2756gat, G2334gat, G2476gat);
nand NAND2_510 (G2757gat, G2331gat, G2477gat);
and AND2_511 (G2758gat, G1520gat, G2481gat);
and AND2_512 (G2761gat, G1722gat, G2482gat);
and AND2_513 (G2764gat, G2478gat, G1770gat);
or OR3_514 (G2768gat, G2486gat, G1789gat, G1790gat);
or OR3_515 (G2769gat, G2487gat, G1797gat, G1798gat);
and AND2_516 (G2898gat, G665gat, G2633gat);
and AND2_517 (G2899gat, G679gat, G2635gat);
and AND2_518 (G2900gat, G686gat, G2637gat);
and AND2_519 (G2901gat, G702gat, G2639gat);
not NOT1_520 (G2962gat, G2746gat);
nand NAND2_521 (G2966gat, G2748gat, G2749gat);
nand NAND2_522 (G2967gat, G2750gat, G2751gat);
nand NAND2_523 (G2973gat, G2754gat, G2755gat);
nand NAND2_524 (G2977gat, G2756gat, G2757gat);
and AND2_525 (G2980gat, G2471gat, G2143gat);
not NOT1_526 (G2984gat, G2488gat);
not NOT1_527 (G2985gat, G2497gat);
not NOT1_528 (G2986gat, G2506gat);
not NOT1_529 (G2987gat, G2515gat);
not NOT1_530 (G2988gat, G2524gat);
not NOT1_531 (G2989gat, G2533gat);
not NOT1_532 (G2990gat, G2542gat);
not NOT1_533 (G2991gat, G2551gat);
not NOT1_534 (G2992gat, G2488gat);
not NOT1_535 (G2993gat, G2497gat);
not NOT1_536 (G2994gat, G2506gat);
not NOT1_537 (G2995gat, G2515gat);
not NOT1_538 (G2996gat, G2524gat);
not NOT1_539 (G2997gat, G2533gat);
not NOT1_540 (G2998gat, G2542gat);
not NOT1_541 (G2999gat, G2551gat);
not NOT1_542 (G3000gat, G2488gat);
not NOT1_543 (G3001gat, G2497gat);
not NOT1_544 (G3002gat, G2506gat);
not NOT1_545 (G3003gat, G2515gat);
not NOT1_546 (G3004gat, G2524gat);
not NOT1_547 (G3005gat, G2533gat);
not NOT1_548 (G3006gat, G2542gat);
not NOT1_549 (G3007gat, G2551gat);
not NOT1_550 (G3008gat, G2488gat);
not NOT1_551 (G3009gat, G2497gat);
not NOT1_552 (G3010gat, G2506gat);
not NOT1_553 (G3011gat, G2515gat);
not NOT1_554 (G3012gat, G2524gat);
not NOT1_555 (G3013gat, G2533gat);
not NOT1_556 (G3014gat, G2542gat);
not NOT1_557 (G3015gat, G2551gat);
not NOT1_558 (G3016gat, G2488gat);
not NOT1_559 (G3017gat, G2497gat);
not NOT1_560 (G3018gat, G2506gat);
not NOT1_561 (G3019gat, G2515gat);
not NOT1_562 (G3020gat, G2524gat);
not NOT1_563 (G3021gat, G2533gat);
not NOT1_564 (G3022gat, G2542gat);
not NOT1_565 (G3023gat, G2551gat);
not NOT1_566 (G3024gat, G2488gat);
not NOT1_567 (G3025gat, G2497gat);
not NOT1_568 (G3026gat, G2506gat);
not NOT1_569 (G3027gat, G2515gat);
not NOT1_570 (G3028gat, G2524gat);
not NOT1_571 (G3029gat, G2533gat);
not NOT1_572 (G3030gat, G2542gat);
not NOT1_573 (G3031gat, G2551gat);
not NOT1_574 (G3032gat, G2488gat);
not NOT1_575 (G3033gat, G2497gat);
not NOT1_576 (G3034gat, G2506gat);
not NOT1_577 (G3035gat, G2515gat);
not NOT1_578 (G3036gat, G2524gat);
not NOT1_579 (G3037gat, G2533gat);
not NOT1_580 (G3038gat, G2542gat);
not NOT1_581 (G3039gat, G2551gat);
not NOT1_582 (G3040gat, G2488gat);
not NOT1_583 (G3041gat, G2497gat);
not NOT1_584 (G3042gat, G2506gat);
not NOT1_585 (G3043gat, G2515gat);
not NOT1_586 (G3044gat, G2524gat);
not NOT1_587 (G3045gat, G2533gat);
not NOT1_588 (G3046gat, G2542gat);
not NOT1_589 (G3047gat, G2551gat);
not NOT1_590 (G3048gat, G2560gat);
not NOT1_591 (G3049gat, G2569gat);
not NOT1_592 (G3050gat, G2578gat);
not NOT1_593 (G3051gat, G2587gat);
not NOT1_594 (G3052gat, G2596gat);
not NOT1_595 (G3053gat, G2605gat);
not NOT1_596 (G3054gat, G2614gat);
not NOT1_597 (G3055gat, G2623gat);
not NOT1_598 (G3056gat, G2560gat);
not NOT1_599 (G3057gat, G2569gat);
not NOT1_600 (G3058gat, G2578gat);
not NOT1_601 (G3059gat, G2587gat);
not NOT1_602 (G3060gat, G2596gat);
not NOT1_603 (G3061gat, G2605gat);
not NOT1_604 (G3062gat, G2614gat);
not NOT1_605 (G3063gat, G2623gat);
not NOT1_606 (G3064gat, G2560gat);
not NOT1_607 (G3065gat, G2569gat);
not NOT1_608 (G3066gat, G2578gat);
not NOT1_609 (G3067gat, G2587gat);
not NOT1_610 (G3068gat, G2596gat);
not NOT1_611 (G3069gat, G2605gat);
not NOT1_612 (G3070gat, G2614gat);
not NOT1_613 (G3071gat, G2623gat);
not NOT1_614 (G3072gat, G2560gat);
not NOT1_615 (G3073gat, G2569gat);
not NOT1_616 (G3074gat, G2578gat);
not NOT1_617 (G3075gat, G2587gat);
not NOT1_618 (G3076gat, G2596gat);
not NOT1_619 (G3077gat, G2605gat);
not NOT1_620 (G3078gat, G2614gat);
not NOT1_621 (G3079gat, G2623gat);
not NOT1_622 (G3080gat, G2560gat);
not NOT1_623 (G3081gat, G2569gat);
not NOT1_624 (G3082gat, G2578gat);
not NOT1_625 (G3083gat, G2587gat);
not NOT1_626 (G3084gat, G2596gat);
not NOT1_627 (G3085gat, G2605gat);
not NOT1_628 (G3086gat, G2614gat);
not NOT1_629 (G3087gat, G2623gat);
not NOT1_630 (G3088gat, G2560gat);
not NOT1_631 (G3089gat, G2569gat);
not NOT1_632 (G3090gat, G2578gat);
not NOT1_633 (G3091gat, G2587gat);
not NOT1_634 (G3092gat, G2596gat);
not NOT1_635 (G3093gat, G2605gat);
not NOT1_636 (G3094gat, G2614gat);
not NOT1_637 (G3095gat, G2623gat);
not NOT1_638 (G3096gat, G2560gat);
not NOT1_639 (G3097gat, G2569gat);
not NOT1_640 (G3098gat, G2578gat);
not NOT1_641 (G3099gat, G2587gat);
not NOT1_642 (G3100gat, G2596gat);
not NOT1_643 (G3101gat, G2605gat);
not NOT1_644 (G3102gat, G2614gat);
not NOT1_645 (G3103gat, G2623gat);
not NOT1_646 (G3104gat, G2560gat);
not NOT1_647 (G3105gat, G2569gat);
not NOT1_648 (G3106gat, G2578gat);
not NOT1_649 (G3107gat, G2587gat);
not NOT1_650 (G3108gat, G2596gat);
not NOT1_651 (G3109gat, G2605gat);
not NOT1_652 (G3110gat, G2614gat);
not NOT1_653 (G3111gat, G2623gat);
not NOT1_654 (G3115gat, G2656gat);
not NOT1_655 (G3118gat, G2652gat);
and AND2_656 (G3119gat, G2768gat, G1674gat);
not NOT1_657 (G3125gat, G2659gat);
not NOT1_658 (G3131gat, G2670gat);
not NOT1_659 (G3134gat, G2666gat);
not NOT1_660 (G3138gat, G2681gat);
not NOT1_661 (G3141gat, G2677gat);
not NOT1_662 (G3145gat, G2692gat);
not NOT1_663 (G3148gat, G2688gat);
and AND2_664 (G3149gat, G2769gat, G1678gat);
not NOT1_665 (G3155gat, G2697gat);
not NOT1_666 (G3161gat, G2710gat);
not NOT1_667 (G3164gat, G2706gat);
not NOT1_668 (G3168gat, G2723gat);
not NOT1_669 (G3171gat, G2719gat);
and AND2_670 (G3172gat, G1909gat, G2648gat);
and AND2_671 (G3175gat, G1913gat, G2662gat);
and AND2_672 (G3178gat, G1913gat, G2673gat);
and AND2_673 (G3181gat, G1913gat, G2684gat);
and AND2_674 (G3184gat, G1922gat, G2702gat);
and AND2_675 (G3187gat, G1922gat, G2715gat);
not NOT1_676 (G3190gat, G2692gat);
not NOT1_677 (G3191gat, G2697gat);
not NOT1_678 (G3192gat, G2710gat);
not NOT1_679 (G3193gat, G2723gat);
and AND5_680 (G3194gat, G2692gat, G2697gat, G2710gat, G2723gat, G1459gat);
nand NAND2_681 (G3195gat, G2745gat, G2962gat);
not NOT1_682 (G3196gat, G2966gat);
or OR3_683 (G3206gat, G2980gat, G2145gat, G2347gat);
and AND2_684 (G3207gat, G124gat, G2984gat);
and AND2_685 (G3208gat, G159gat, G2985gat);
and AND2_686 (G3209gat, G150gat, G2986gat);
and AND2_687 (G3210gat, G143gat, G2987gat);
and AND2_688 (G3211gat, G137gat, G2988gat);
and AND2_689 (G3212gat, G132gat, G2989gat);
and AND2_690 (G3213gat, G128gat, G2990gat);
and AND2_691 (G3214gat, G125gat, G2991gat);
and AND2_692 (G3215gat, G125gat, G2992gat);
and AND2_693 (G3216gat, G655gat, G2993gat);
and AND2_694 (G3217gat, G159gat, G2994gat);
and AND2_695 (G3218gat, G150gat, G2995gat);
and AND2_696 (G3219gat, G143gat, G2996gat);
and AND2_697 (G3220gat, G137gat, G2997gat);
and AND2_698 (G3221gat, G132gat, G2998gat);
and AND2_699 (G3222gat, G128gat, G2999gat);
and AND2_700 (G3223gat, G128gat, G3000gat);
and AND2_701 (G3224gat, G670gat, G3001gat);
and AND2_702 (G3225gat, G655gat, G3002gat);
and AND2_703 (G3226gat, G159gat, G3003gat);
and AND2_704 (G3227gat, G150gat, G3004gat);
and AND2_705 (G3228gat, G143gat, G3005gat);
and AND2_706 (G3229gat, G137gat, G3006gat);
and AND2_707 (G3230gat, G132gat, G3007gat);
and AND2_708 (G3231gat, G132gat, G3008gat);
and AND2_709 (G3232gat, G690gat, G3009gat);
and AND2_710 (G3233gat, G670gat, G3010gat);
and AND2_711 (G3234gat, G655gat, G3011gat);
and AND2_712 (G3235gat, G159gat, G3012gat);
and AND2_713 (G3236gat, G150gat, G3013gat);
and AND2_714 (G3237gat, G143gat, G3014gat);
and AND2_715 (G3238gat, G137gat, G3015gat);
and AND2_716 (G3239gat, G137gat, G3016gat);
and AND2_717 (G3240gat, G706gat, G3017gat);
and AND2_718 (G3241gat, G690gat, G3018gat);
and AND2_719 (G3242gat, G670gat, G3019gat);
and AND2_720 (G3243gat, G655gat, G3020gat);
and AND2_721 (G3244gat, G159gat, G3021gat);
and AND2_722 (G3245gat, G150gat, G3022gat);
and AND2_723 (G3246gat, G143gat, G3023gat);
and AND2_724 (G3247gat, G143gat, G3024gat);
and AND2_725 (G3248gat, G715gat, G3025gat);
and AND2_726 (G3249gat, G706gat, G3026gat);
and AND2_727 (G3250gat, G690gat, G3027gat);
and AND2_728 (G3251gat, G670gat, G3028gat);
and AND2_729 (G3252gat, G655gat, G3029gat);
and AND2_730 (G3253gat, G159gat, G3030gat);
and AND2_731 (G3254gat, G150gat, G3031gat);
and AND2_732 (G3255gat, G150gat, G3032gat);
and AND2_733 (G3256gat, G727gat, G3033gat);
and AND2_734 (G3257gat, G715gat, G3034gat);
and AND2_735 (G3258gat, G706gat, G3035gat);
and AND2_736 (G3259gat, G690gat, G3036gat);
and AND2_737 (G3260gat, G670gat, G3037gat);
and AND2_738 (G3261gat, G655gat, G3038gat);
and AND2_739 (G3262gat, G159gat, G3039gat);
and AND2_740 (G3263gat, G159gat, G3040gat);
and AND2_741 (G3264gat, G740gat, G3041gat);
and AND2_742 (G3265gat, G727gat, G3042gat);
and AND2_743 (G3266gat, G715gat, G3043gat);
and AND2_744 (G3267gat, G706gat, G3044gat);
and AND2_745 (G3268gat, G690gat, G3045gat);
and AND2_746 (G3269gat, G670gat, G3046gat);
and AND2_747 (G3270gat, G655gat, G3047gat);
and AND2_748 (G3271gat, G283gat, G3048gat);
and AND2_749 (G3272gat, G670gat, G3049gat);
and AND2_750 (G3273gat, G690gat, G3050gat);
and AND2_751 (G3274gat, G706gat, G3051gat);
and AND2_752 (G3275gat, G715gat, G3052gat);
and AND2_753 (G3276gat, G727gat, G3053gat);
and AND2_754 (G3277gat, G740gat, G3054gat);
and AND2_755 (G3278gat, G753gat, G3055gat);
and AND2_756 (G3279gat, G294gat, G3056gat);
and AND2_757 (G3280gat, G690gat, G3057gat);
and AND2_758 (G3281gat, G706gat, G3058gat);
and AND2_759 (G3282gat, G715gat, G3059gat);
and AND2_760 (G3283gat, G727gat, G3060gat);
and AND2_761 (G3284gat, G740gat, G3061gat);
and AND2_762 (G3285gat, G753gat, G3062gat);
and AND2_763 (G3286gat, G283gat, G3063gat);
and AND2_764 (G3287gat, G303gat, G3064gat);
and AND2_765 (G3288gat, G706gat, G3065gat);
and AND2_766 (G3289gat, G715gat, G3066gat);
and AND2_767 (G3290gat, G727gat, G3067gat);
and AND2_768 (G3291gat, G740gat, G3068gat);
and AND2_769 (G3292gat, G753gat, G3069gat);
and AND2_770 (G3293gat, G283gat, G3070gat);
and AND2_771 (G3294gat, G294gat, G3071gat);
and AND2_772 (G3295gat, G311gat, G3072gat);
and AND2_773 (G3296gat, G715gat, G3073gat);
and AND2_774 (G3297gat, G727gat, G3074gat);
and AND2_775 (G3298gat, G740gat, G3075gat);
and AND2_776 (G3299gat, G753gat, G3076gat);
and AND2_777 (G3300gat, G283gat, G3077gat);
and AND2_778 (G3301gat, G294gat, G3078gat);
and AND2_779 (G3302gat, G303gat, G3079gat);
and AND2_780 (G3303gat, G317gat, G3080gat);
and AND2_781 (G3304gat, G727gat, G3081gat);
and AND2_782 (G3305gat, G740gat, G3082gat);
and AND2_783 (G3306gat, G753gat, G3083gat);
and AND2_784 (G3307gat, G283gat, G3084gat);
and AND2_785 (G3308gat, G294gat, G3085gat);
and AND2_786 (G3309gat, G303gat, G3086gat);
and AND2_787 (G3310gat, G311gat, G3087gat);
and AND2_788 (G3311gat, G322gat, G3088gat);
and AND2_789 (G3312gat, G740gat, G3089gat);
and AND2_790 (G3313gat, G753gat, G3090gat);
and AND2_791 (G3314gat, G283gat, G3091gat);
and AND2_792 (G3315gat, G294gat, G3092gat);
and AND2_793 (G3316gat, G303gat, G3093gat);
and AND2_794 (G3317gat, G311gat, G3094gat);
and AND2_795 (G3318gat, G317gat, G3095gat);
and AND2_796 (G3319gat, G326gat, G3096gat);
and AND2_797 (G3320gat, G753gat, G3097gat);
and AND2_798 (G3321gat, G283gat, G3098gat);
and AND2_799 (G3322gat, G294gat, G3099gat);
and AND2_800 (G3323gat, G303gat, G3100gat);
and AND2_801 (G3324gat, G311gat, G3101gat);
and AND2_802 (G3325gat, G317gat, G3102gat);
and AND2_803 (G3326gat, G322gat, G3103gat);
and AND2_804 (G3327gat, G329gat, G3104gat);
and AND2_805 (G3328gat, G283gat, G3105gat);
and AND2_806 (G3329gat, G294gat, G3106gat);
and AND2_807 (G3330gat, G303gat, G3107gat);
and AND2_808 (G3331gat, G311gat, G3108gat);
and AND2_809 (G3332gat, G317gat, G3109gat);
and AND2_810 (G3333gat, G322gat, G3110gat);
and AND2_811 (G3334gat, G326gat, G3111gat);
and AND5_812 (G3383gat, G3190gat, G3191gat, G3192gat, G3193gat, G917gat);
and AND2_813 (G3387gat, G3196gat, G1736gat);
and AND2_814 (G3388gat, G2977gat, G2149gat);
and AND2_815 (G3389gat, G2973gat, G1737gat);
or OR4_816 (G33890gat, G3207gat, G3208gat, G3209gat, G3210gat);
or OR4_817 (G33891gat, G3211gat, G3212gat, G3213gat, G3214gat);
nor NOR2_818 (G3390gat, G33890gat, G33891gat);
or OR4_819 (G33900gat, G3215gat, G3216gat, G3217gat, G3218gat);
or OR4_820 (G33901gat, G3219gat, G3220gat, G3221gat, G3222gat);
nor NOR2_821 (G3391gat, G33900gat, G33901gat);
or OR4_822 (G33910gat, G3223gat, G3224gat, G3225gat, G3226gat);
or OR4_823 (G33911gat, G3227gat, G3228gat, G3229gat, G3230gat);
nor NOR2_824 (G3392gat, G33910gat, G33911gat);
or OR4_825 (G33920gat, G3231gat, G3232gat, G3233gat, G3234gat);
or OR4_826 (G33921gat, G3235gat, G3236gat, G3237gat, G3238gat);
nor NOR2_827 (G3393gat, G33920gat, G33921gat);
or OR4_828 (G33930gat, G3239gat, G3240gat, G3241gat, G3242gat);
or OR4_829 (G33931gat, G3243gat, G3244gat, G3245gat, G3246gat);
nor NOR2_830 (G3394gat, G33930gat, G33931gat);
or OR4_831 (G33940gat, G3247gat, G3248gat, G3249gat, G3250gat);
or OR4_832 (G33941gat, G3251gat, G3252gat, G3253gat, G3254gat);
nor NOR2_833 (G3395gat, G33940gat, G33941gat);
or OR4_834 (G33950gat, G3255gat, G3256gat, G3257gat, G3258gat);
or OR4_835 (G33951gat, G3259gat, G3260gat, G3261gat, G3262gat);
nor NOR2_836 (G3396gat, G33950gat, G33951gat);
or OR4_837 (G33960gat, G3263gat, G3264gat, G3265gat, G3266gat);
or OR4_838 (G33961gat, G3267gat, G3268gat, G3269gat, G3270gat);
nor NOR2_839 (G3397gat, G33960gat, G33961gat);
or OR4_840 (G33970gat, G3271gat, G3272gat, G3273gat, G3274gat);
or OR4_841 (G33971gat, G3275gat, G3276gat, G3277gat, G3278gat);
nor NOR2_842 (G3398gat, G33970gat, G33971gat);
or OR4_843 (G33980gat, G3279gat, G3280gat, G3281gat, G3282gat);
or OR4_844 (G33981gat, G3283gat, G3284gat, G3285gat, G3286gat);
nor NOR2_845 (G3399gat, G33980gat, G33981gat);
or OR4_846 (G33990gat, G3287gat, G3288gat, G3289gat, G3290gat);
or OR4_847 (G33991gat, G3291gat, G3292gat, G3293gat, G3294gat);
nor NOR2_848 (G3400gat, G33990gat, G33991gat);
or OR4_849 (G34000gat, G3295gat, G3296gat, G3297gat, G3298gat);
or OR4_850 (G34001gat, G3299gat, G3300gat, G3301gat, G3302gat);
nor NOR2_851 (G3401gat, G34000gat, G34001gat);
or OR4_852 (G34010gat, G3303gat, G3304gat, G3305gat, G3306gat);
or OR4_853 (G34011gat, G3307gat, G3308gat, G3309gat, G3310gat);
nor NOR2_854 (G3402gat, G34010gat, G34011gat);
or OR4_855 (G34020gat, G3311gat, G3312gat, G3313gat, G3314gat);
or OR4_856 (G34021gat, G3315gat, G3316gat, G3317gat, G3318gat);
nor NOR2_857 (G3403gat, G34020gat, G34021gat);
or OR4_858 (G34030gat, G3319gat, G3320gat, G3321gat, G3322gat);
or OR4_859 (G34031gat, G3323gat, G3324gat, G3325gat, G3326gat);
nor NOR2_860 (G3404gat, G34030gat, G34031gat);
or OR4_861 (G34040gat, G3327gat, G3328gat, G3329gat, G3330gat);
or OR4_862 (G34041gat, G3331gat, G3332gat, G3333gat, G3334gat);
nor NOR2_863 (G3405gat, G34040gat, G34041gat);
and AND2_864 (G3406gat, G3206gat, G2641gat);
and AND3_865 (G3407gat, G169gat, G2648gat, G3112gat);
and AND3_866 (G3410gat, G179gat, G2648gat, G3115gat);
and AND3_867 (G3413gat, G190gat, G2652gat, G3115gat);
and AND3_868 (G3414gat, G200gat, G2652gat, G3112gat);
or OR3_869 (G3415gat, G3119gat, G1875gat, G2073gat);
nor NOR3_870 (G3419gat, G3119gat, G1875gat, G2073gat);
and AND3_871 (G3423gat, G169gat, G2662gat, G3128gat);
and AND3_872 (G3426gat, G179gat, G2662gat, G3131gat);
and AND3_873 (G3429gat, G190gat, G2666gat, G3131gat);
and AND3_874 (G3430gat, G200gat, G2666gat, G3128gat);
and AND3_875 (G3431gat, G169gat, G2673gat, G3135gat);
and AND3_876 (G3434gat, G179gat, G2673gat, G3138gat);
and AND3_877 (G3437gat, G190gat, G2677gat, G3138gat);
and AND3_878 (G3438gat, G200gat, G2677gat, G3135gat);
and AND3_879 (G3439gat, G169gat, G2684gat, G3142gat);
and AND3_880 (G3442gat, G179gat, G2684gat, G3145gat);
and AND3_881 (G3445gat, G190gat, G2688gat, G3145gat);
and AND3_882 (G3446gat, G200gat, G2688gat, G3142gat);
or OR3_883 (G3447gat, G3149gat, G1895gat, G2093gat);
nor NOR3_884 (G3451gat, G3149gat, G1895gat, G2093gat);
and AND3_885 (G3455gat, G169gat, G2702gat, G3158gat);
and AND3_886 (G3458gat, G179gat, G2702gat, G3161gat);
and AND3_887 (G3461gat, G190gat, G2706gat, G3161gat);
and AND3_888 (G3462gat, G200gat, G2706gat, G3158gat);
and AND3_889 (G3463gat, G169gat, G2715gat, G3165gat);
and AND3_890 (G3466gat, G179gat, G2715gat, G3168gat);
and AND3_891 (G3469gat, G190gat, G2719gat, G3168gat);
and AND3_892 (G3470gat, G200gat, G2719gat, G3165gat);
or OR2_893 (G3471gat, G3194gat, G3383gat);
nor NOR2_894 (G3534gat, G3387gat, G2350gat);
or OR3_895 (G3535gat, G3388gat, G2151gat, G2351gat);
nor NOR2_896 (G3536gat, G3389gat, G1966gat);
and AND2_897 (G3537gat, G3390gat, G2209gat);
and AND2_898 (G3538gat, G3398gat, G2210gat);
and AND2_899 (G3539gat, G3391gat, G1842gat);
and AND2_900 (G3540gat, G3399gat, G1369gat);
and AND2_901 (G3541gat, G3392gat, G1843gat);
and AND2_902 (G3542gat, G3400gat, G1369gat);
and AND2_903 (G3543gat, G3393gat, G1844gat);
and AND2_904 (G3544gat, G3401gat, G1369gat);
and AND2_905 (G3545gat, G3394gat, G1845gat);
and AND2_906 (G3546gat, G3402gat, G1369gat);
and AND2_907 (G3547gat, G3395gat, G1846gat);
and AND2_908 (G3548gat, G3403gat, G1369gat);
and AND2_909 (G3549gat, G3396gat, G1847gat);
and AND2_910 (G3550gat, G3404gat, G1369gat);
and AND2_911 (G3551gat, G3397gat, G1848gat);
and AND2_912 (G3552gat, G3405gat, G1369gat);
or OR3_913 (G3557gat, G3413gat, G3414gat, G3118gat);
or OR3_914 (G3568gat, G3429gat, G3430gat, G3134gat);
or OR3_915 (G3573gat, G3437gat, G3438gat, G3141gat);
or OR3_916 (G3578gat, G3445gat, G3446gat, G3148gat);
or OR3_917 (G3589gat, G3461gat, G3462gat, G3164gat);
or OR3_918 (G3594gat, G3469gat, G3470gat, G3171gat);
and AND2_919 (G3605gat, G3471gat, G2728gat);
not NOT1_920 (G3626gat, G3478gat);
not NOT1_921 (G3627gat, G3481gat);
not NOT1_922 (G3628gat, G3487gat);
not NOT1_923 (G3629gat, G3484gat);
not NOT1_924 (G3630gat, G3472gat);
not NOT1_925 (G3631gat, G3475gat);
and AND2_926 (G3632gat, G3536gat, G2152gat);
and AND2_927 (G3633gat, G3534gat, G2155gat);
or OR3_928 (G3634gat, G3537gat, G3538gat, G2398gat);
or OR2_929 (G3635gat, G3539gat, G3540gat);
or OR2_930 (G3636gat, G3541gat, G3542gat);
or OR2_931 (G3637gat, G3543gat, G3544gat);
or OR2_932 (G3638gat, G3545gat, G3546gat);
or OR2_933 (G3639gat, G3547gat, G3548gat);
or OR2_934 (G3640gat, G3549gat, G3550gat);
or OR2_935 (G3641gat, G3551gat, G3552gat);
and AND2_936 (G3642gat, G3535gat, G2643gat);
or OR2_937 (G3643gat, G3407gat, G3410gat);
nor NOR2_938 (G3644gat, G3407gat, G3410gat);
and AND3_939 (G3645gat, G169gat, G3415gat, G3122gat);
and AND3_940 (G3648gat, G179gat, G3415gat, G3125gat);
and AND3_941 (G3651gat, G190gat, G3419gat, G3125gat);
and AND3_942 (G3652gat, G200gat, G3419gat, G3122gat);
not NOT1_943 (G3653gat, G3419gat);
or OR2_944 (G3654gat, G3423gat, G3426gat);
nor NOR2_945 (G3657gat, G3423gat, G3426gat);
or OR2_946 (G3658gat, G3431gat, G3434gat);
nor NOR2_947 (G3661gat, G3431gat, G3434gat);
or OR2_948 (G3662gat, G3439gat, G3442gat);
nor NOR2_949 (G3663gat, G3439gat, G3442gat);
and AND3_950 (G3664gat, G169gat, G3447gat, G3152gat);
and AND3_951 (G3667gat, G179gat, G3447gat, G3155gat);
and AND3_952 (G3670gat, G190gat, G3451gat, G3155gat);
and AND3_953 (G3671gat, G200gat, G3451gat, G3152gat);
not NOT1_954 (G3672gat, G3451gat);
or OR2_955 (G3673gat, G3455gat, G3458gat);
nor NOR2_956 (G3676gat, G3455gat, G3458gat);
or OR2_957 (G3677gat, G3463gat, G3466gat);
nor NOR2_958 (G3680gat, G3463gat, G3466gat);
not NOT1_959 (G3681gat, G3493gat);
and AND2_960 (G3682gat, G1909gat, G3415gat);
not NOT1_961 (G3685gat, G3496gat);
not NOT1_962 (G3686gat, G3499gat);
not NOT1_963 (G3687gat, G3502gat);
not NOT1_964 (G3688gat, G3505gat);
not NOT1_965 (G3689gat, G3511gat);
and AND2_966 (G3690gat, G1922gat, G3447gat);
not NOT1_967 (G3693gat, G3517gat);
not NOT1_968 (G3694gat, G3520gat);
not NOT1_969 (G3695gat, G3523gat);
not NOT1_970 (G3696gat, G3514gat);
not NOT1_971 (G3703gat, G3490gat);
not NOT1_972 (G3704gat, G3508gat);
nand NAND2_973 (G3705gat, G3475gat, G3630gat);
nand NAND2_974 (G3706gat, G3472gat, G3631gat);
nand NAND2_975 (G3707gat, G3481gat, G3626gat);
nand NAND2_976 (G3708gat, G3478gat, G3627gat);
or OR3_977 (G3711gat, G3632gat, G2352gat, G2353gat);
or OR3_978 (G3712gat, G3633gat, G2354gat, G2355gat);
and AND2_979 (G3713gat, G3634gat, G2632gat);
and AND2_980 (G3714gat, G3635gat, G2634gat);
and AND2_981 (G3715gat, G3636gat, G2636gat);
and AND2_982 (G3716gat, G3637gat, G2638gat);
and AND2_983 (G3717gat, G3638gat, G2640gat);
and AND2_984 (G3718gat, G3639gat, G2642gat);
and AND2_985 (G3719gat, G3640gat, G2644gat);
and AND2_986 (G3720gat, G3641gat, G2646gat);
and AND2_987 (G3721gat, G3644gat, G3557gat);
or OR3_988 (G3731gat, G3651gat, G3652gat, G3653gat);
and AND2_989 (G3734gat, G3657gat, G3568gat);
and AND2_990 (G3740gat, G3661gat, G3573gat);
and AND2_991 (G3743gat, G3663gat, G3578gat);
or OR3_992 (G3753gat, G3670gat, G3671gat, G3672gat);
and AND2_993 (G3756gat, G3676gat, G3589gat);
and AND2_994 (G3762gat, G3680gat, G3594gat);
not NOT1_995 (G3765gat, G3643gat);
not NOT1_996 (G3766gat, G3662gat);
nand NAND2_997 (G3773gat, G3705gat, G3706gat);
nand NAND2_998 (G3774gat, G3707gat, G3708gat);
nand NAND2_999 (G3775gat, G3700gat, G3628gat);
not NOT1_1000 (G3776gat, G3700gat);
nand NAND2_1001 (G3777gat, G3697gat, G3629gat);
not NOT1_1002 (G3778gat, G3697gat);
and AND2_1003 (G3779gat, G3712gat, G2645gat);
and AND2_1004 (G3780gat, G3711gat, G2647gat);
or OR2_1005 (G3786gat, G3645gat, G3648gat);
nor NOR2_1006 (G3789gat, G3645gat, G3648gat);
or OR2_1007 (G3800gat, G3664gat, G3667gat);
nor NOR2_1008 (G3803gat, G3664gat, G3667gat);
and AND2_1009 (G3809gat, G3654gat, G1917gat);
and AND2_1010 (G3812gat, G3658gat, G1917gat);
and AND2_1011 (G3815gat, G3673gat, G1926gat);
and AND2_1012 (G3818gat, G3677gat, G1926gat);
nand NAND2_1013 (G3833gat, G3773gat, G3774gat);
nand NAND2_1014 (G3834gat, G3487gat, G3776gat);
nand NAND2_1015 (G3835gat, G3484gat, G3778gat);
and AND2_1016 (G3838gat, G3789gat, G3731gat);
and AND2_1017 (G3845gat, G3803gat, G3753gat);
nand NAND2_1018 (G3884gat, G3775gat, G3834gat);
nand NAND2_1019 (G3885gat, G3777gat, G3835gat);
nand NAND2_1020 (G3894gat, G3721gat, G3786gat);
nand NAND2_1021 (G3895gat, G3743gat, G3800gat);
not NOT1_1022 (G3898gat, G3821gat);
not NOT1_1023 (G3899gat, G3824gat);
not NOT1_1024 (G3906gat, G3830gat);
not NOT1_1025 (G3911gat, G3827gat);
and AND2_1026 (G3912gat, G3786gat, G1912gat);
and AND2_1027 (G3916gat, G3800gat, G1917gat);
not NOT1_1028 (G3920gat, G3809gat);
not NOT1_1029 (G3924gat, G3884gat);
not NOT1_1030 (G3925gat, G3885gat);
and AND4_1031 (G3926gat, G3721gat, G3838gat, G3734gat, G3740gat);
nand NAND3_1032 (G3930gat, G3721gat, G3838gat, G3654gat);
nand NAND4_1033 (G3931gat, G3658gat, G3838gat, G3734gat, G3721gat);
and AND4_1034 (G3932gat, G3743gat, G3845gat, G3756gat, G3762gat);
nand NAND3_1035 (G3935gat, G3743gat, G3845gat, G3673gat);
nand NAND4_1036 (G3936gat, G3677gat, G3845gat, G3756gat, G3743gat);
not NOT1_1037 (G3947gat, G3912gat);
not NOT1_1038 (G3948gat, G3916gat);
nand NAND2_1039 (G3987gat, G3924gat, G3925gat);
nand NAND4_1040 (G3992gat, G3765gat, G3894gat, G3930gat, G3931gat);
nand NAND4_1041 (G3996gat, G3766gat, G3895gat, G3935gat, G3936gat);
not NOT1_1042 (G4013gat, G3921gat);
and AND2_1043 (G4028gat, G3932gat, G3926gat);
nand NAND2_1044 (G4029gat, G3953gat, G3681gat);
nand NAND2_1045 (G4030gat, G3959gat, G3686gat);
nand NAND2_1046 (G4031gat, G3965gat, G3688gat);
nand NAND2_1047 (G4032gat, G3971gat, G3689gat);
nand NAND2_1048 (G4033gat, G3977gat, G3693gat);
nand NAND2_1049 (G4034gat, G3983gat, G3695gat);
not NOT1_1050 (G4042gat, G3953gat);
not NOT1_1051 (G4043gat, G3956gat);
nand NAND2_1052 (G4044gat, G3956gat, G3685gat);
not NOT1_1053 (G4045gat, G3959gat);
not NOT1_1054 (G4046gat, G3962gat);
nand NAND2_1055 (G4047gat, G3962gat, G3687gat);
not NOT1_1056 (G4048gat, G3965gat);
not NOT1_1057 (G4049gat, G3971gat);
not NOT1_1058 (G4050gat, G3977gat);
not NOT1_1059 (G4051gat, G3980gat);
nand NAND2_1060 (G4052gat, G3980gat, G3694gat);
not NOT1_1061 (G4053gat, G3983gat);
not NOT1_1062 (G4054gat, G3974gat);
nand NAND2_1063 (G4055gat, G3974gat, G3696gat);
and AND2_1064 (G4056gat, G3932gat, G2304gat);
not NOT1_1065 (G4057gat, G3950gat);
nand NAND2_1066 (G4058gat, G3950gat, G3703gat);
not NOT1_1067 (G4065gat, G3968gat);
nand NAND2_1068 (G4066gat, G3968gat, G3704gat);
nand NAND2_1069 (G4073gat, G3926gat, G3996gat);
not NOT1_1070 (G4074gat, G3992gat);
nand NAND2_1071 (G4075gat, G3493gat, G4042gat);
nand NAND2_1072 (G4076gat, G3499gat, G4045gat);
nand NAND2_1073 (G4077gat, G3505gat, G4048gat);
nand NAND2_1074 (G4078gat, G3511gat, G4049gat);
nand NAND2_1075 (G4079gat, G3517gat, G4050gat);
nand NAND2_1076 (G4080gat, G3523gat, G4053gat);
nand NAND2_1077 (G4085gat, G3496gat, G4043gat);
nand NAND2_1078 (G4086gat, G3502gat, G4046gat);
nand NAND2_1079 (G4088gat, G3520gat, G4051gat);
nand NAND2_1080 (G4090gat, G3514gat, G4054gat);
and AND2_1081 (G4091gat, G3996gat, G1926gat);
or OR2_1082 (G4094gat, G3605gat, G4056gat);
nand NAND2_1083 (G4098gat, G3490gat, G4057gat);
nand NAND2_1084 (G4101gat, G3508gat, G4065gat);
and AND2_1085 (G4104gat, G4073gat, G4074gat);
nand NAND2_1086 (G4105gat, G4075gat, G4029gat);
nand NAND2_1087 (G4106gat, G4062gat, G3899gat);
nand NAND2_1088 (G4107gat, G4076gat, G4030gat);
nand NAND2_1089 (G4108gat, G4077gat, G4031gat);
nand NAND2_1090 (G4109gat, G4078gat, G4032gat);
nand NAND2_1091 (G4110gat, G4070gat, G3906gat);
nand NAND2_1092 (G4111gat, G4079gat, G4033gat);
nand NAND2_1093 (G4112gat, G4080gat, G4034gat);
not NOT1_1094 (G4113gat, G4059gat);
nand NAND2_1095 (G4114gat, G4059gat, G3898gat);
not NOT1_1096 (G4115gat, G4062gat);
nand NAND2_1097 (G4116gat, G4085gat, G4044gat);
nand NAND2_1098 (G4119gat, G4086gat, G4047gat);
not NOT1_1099 (G4122gat, G4070gat);
nand NAND2_1100 (G4123gat, G4088gat, G4052gat);
not NOT1_1101 (G4126gat, G4067gat);
nand NAND2_1102 (G4127gat, G4067gat, G3911gat);
nand NAND2_1103 (G4128gat, G4090gat, G4055gat);
nand NAND2_1104 (G4139gat, G4098gat, G4058gat);
nand NAND2_1105 (G4142gat, G4101gat, G4066gat);
not NOT1_1106 (G4145gat, G4104gat);
not NOT1_1107 (G4146gat, G4105gat);
nand NAND2_1108 (G4147gat, G3824gat, G4115gat);
not NOT1_1109 (G4148gat, G4107gat);
not NOT1_1110 (G4149gat, G4108gat);
not NOT1_1111 (G4150gat, G4109gat);
nand NAND2_1112 (G4151gat, G3830gat, G4122gat);
not NOT1_1113 (G4152gat, G4111gat);
not NOT1_1114 (G4153gat, G4112gat);
nand NAND2_1115 (G4154gat, G3821gat, G4113gat);
nand NAND2_1116 (G4161gat, G3827gat, G4126gat);
and AND2_1117 (G4186gat, G330gat, G4094gat);
and AND2_1118 (G4189gat, G4146gat, G2230gat);
nand NAND2_1119 (G4190gat, G4147gat, G4106gat);
and AND2_1120 (G4191gat, G4148gat, G2232gat);
and AND2_1121 (G4192gat, G4149gat, G2233gat);
and AND2_1122 (G4193gat, G4150gat, G2234gat);
nand NAND2_1123 (G4194gat, G4151gat, G4110gat);
and AND2_1124 (G4195gat, G4152gat, G2236gat);
and AND2_1125 (G4196gat, G4153gat, G2237gat);
nand NAND2_1126 (G4197gat, G4154gat, G4114gat);
nand NAND2_1127 (G4218gat, G4161gat, G4127gat);
and AND2_1128 (G4238gat, G4128gat, G3917gat);
not NOT1_1129 (G4239gat, G4139gat);
not NOT1_1130 (G4241gat, G4142gat);
and AND2_1131 (G4242gat, G330gat, G4123gat);
nor NOR3_1132 (G4251gat, G3713gat, G4189gat, G2898gat);
not NOT1_1133 (G4252gat, G4190gat);
nor NOR3_1134 (G4253gat, G3715gat, G4191gat, G2900gat);
nor NOR3_1135 (G4254gat, G3716gat, G4192gat, G2901gat);
nor NOR3_1136 (G4255gat, G3717gat, G4193gat, G3406gat);
not NOT1_1137 (G4256gat, G4194gat);
nor NOR3_1138 (G4257gat, G3719gat, G4195gat, G3779gat);
nor NOR3_1139 (G4258gat, G3720gat, G4196gat, G3780gat);
and AND2_1140 (G4283gat, G4167gat, G4035gat);
and AND2_1141 (G4284gat, G4174gat, G4035gat);
or OR2_1142 (G4287gat, G3815gat, G4238gat);
not NOT1_1143 (G4291gat, G4186gat);
not NOT1_1144 (G4295gat, G4167gat);
not NOT1_1145 (G4299gat, G4182gat);
and AND2_1146 (G4303gat, G4252gat, G2231gat);
and AND2_1147 (G4304gat, G4256gat, G2235gat);
or OR2_1148 (G4310gat, G3992gat, G4283gat);
and AND3_1149 (G4316gat, G4174gat, G4213gat, G4203gat);
and AND2_1150 (G4317gat, G4174gat, G4209gat);
and AND3_1151 (G4318gat, G4223gat, G4128gat, G4218gat);
and AND2_1152 (G4319gat, G4223gat, G4128gat);
and AND2_1153 (G4322gat, G4167gat, G4209gat);
nand NAND2_1154 (G4325gat, G4203gat, G3913gat);
nand NAND3_1155 (G4326gat, G4203gat, G4213gat, G4167gat);
nand NAND2_1156 (G4327gat, G4218gat, G3815gat);
nand NAND3_1157 (G4328gat, G4218gat, G4128gat, G3917gat);
nand NAND2_1158 (G4329gat, G4247gat, G4013gat);
not NOT1_1159 (G4330gat, G4247gat);
and AND3_1160 (G4331gat, G330gat, G4094gat, G4295gat);
and AND2_1161 (G4335gat, G4251gat, G2730gat);
and AND2_1162 (G4338gat, G4253gat, G2734gat);
and AND2_1163 (G4341gat, G4254gat, G2736gat);
and AND2_1164 (G4344gat, G4255gat, G2738gat);
and AND2_1165 (G4347gat, G4257gat, G2742gat);
and AND2_1166 (G4350gat, G4258gat, G2744gat);
and AND2_1167 (G4371gat, G4223gat, G4223gat);
nor NOR3_1168 (G4376gat, G3714gat, G4303gat, G2899gat);
nor NOR3_1169 (G4377gat, G3718gat, G4304gat, G3642gat);
and AND2_1170 (G4387gat, G330gat, G4317gat);
and AND2_1171 (G4390gat, G330gat, G4318gat);
nand NAND2_1172 (G4393gat, G3921gat, G4330gat);
nand NAND3_1173 (G4416gat, G3920gat, G4325gat, G4326gat);
or OR2_1174 (G4421gat, G3812gat, G4322gat);
nand NAND3_1175 (G4427gat, G3948gat, G4327gat, G4328gat);
and AND2_1176 (G4435gat, G330gat, G4316gat);
or OR2_1177 (G4442gat, G4331gat, G4296gat);
and AND4_1178 (G4443gat, G4174gat, G4305gat, G4203gat, G4213gat);
nand NAND2_1179 (G4446gat, G4305gat, G3809gat);
nand NAND3_1180 (G4447gat, G4305gat, G4200gat, G3913gat);
nand NAND4_1181 (G4448gat, G4305gat, G4200gat, G4213gat, G4167gat);
not NOT1_1182 (G4452gat, G4356gat);
nand NAND2_1183 (G4458gat, G4329gat, G4393gat);
not NOT1_1184 (G4461gat, G4365gat);
not NOT1_1185 (G4462gat, G4368gat);
nand NAND2_1186 (G4463gat, G4371gat, G1460gat);
not NOT1_1187 (G4464gat, G4371gat);
nor NOR2_1188 (G4468gat, G4331gat, G4296gat);
and AND2_1189 (G4472gat, G4376gat, G2732gat);
and AND2_1190 (G4475gat, G4377gat, G2740gat);
not NOT1_1191 (G4484gat, G4353gat);
not NOT1_1192 (G4486gat, G4359gat);
nand NAND2_1193 (G4487gat, G4359gat, G4299gat);
not NOT1_1194 (G4491gat, G4362gat);
and AND2_1195 (G4493gat, G330gat, G4319gat);
not NOT1_1196 (G4496gat, G4398gat);
and AND2_1197 (G4497gat, G4287gat, G4398gat);
and AND2_1198 (G4498gat, G4442gat, G1769gat);
nand NAND4_1199 (G4503gat, G3947gat, G4446gat, G4447gat, G4448gat);
not NOT1_1200 (G4506gat, G4413gat);
not NOT1_1201 (G4507gat, G4435gat);
not NOT1_1202 (G4508gat, G4421gat);
nand NAND2_1203 (G4509gat, G4421gat, G4452gat);
not NOT1_1204 (G4510gat, G4427gat);
nand NAND2_1205 (G4511gat, G4427gat, G4241gat);
nand NAND2_1206 (G4515gat, G965gat, G4464gat);
not NOT1_1207 (G4526gat, G4416gat);
nand NAND2_1208 (G4527gat, G4416gat, G4484gat);
nand NAND2_1209 (G4528gat, G4182gat, G4486gat);
not NOT1_1210 (G4529gat, G4430gat);
nand NAND2_1211 (G4530gat, G4430gat, G4491gat);
and AND3_1212 (G4545gat, G330gat, G4319gat, G4496gat);
and AND2_1213 (G4549gat, G330gat, G4443gat);
nand NAND2_1214 (G4552gat, G4356gat, G4508gat);
nand NAND2_1215 (G4555gat, G4142gat, G4510gat);
not NOT1_1216 (G4558gat, G4493gat);
nand NAND2_1217 (G4559gat, G4463gat, G4515gat);
not NOT1_1218 (G4562gat, G4465gat);
and AND2_1219 (G4563gat, G4310gat, G4465gat);
not NOT1_1220 (G4568gat, G4479gat);
nand NAND2_1221 (G4572gat, G4353gat, G4526gat);
nand NAND2_1222 (G4573gat, G4362gat, G4529gat);
nand NAND2_1223 (G4576gat, G4487gat, G4528gat);
or OR3_1224 (G4587gat, G2758gat, G4498gat, G2761gat);
nor NOR3_1225 (G4588gat, G2758gat, G4498gat, G2761gat);
or OR2_1226 (G4589gat, G4545gat, G4497gat);
nand NAND2_1227 (G4593gat, G4552gat, G4509gat);
not NOT1_1228 (G4596gat, G4531gat);
not NOT1_1229 (G4597gat, G4534gat);
nand NAND2_1230 (G4599gat, G4555gat, G4511gat);
not NOT1_1231 (G4602gat, G4537gat);
not NOT1_1232 (G4603gat, G4540gat);
and AND3_1233 (G4608gat, G330gat, G4284gat, G4562gat);
nand NAND2_1234 (G4619gat, G4572gat, G4527gat);
nand NAND2_1235 (G4623gat, G4573gat, G4530gat);
not NOT1_1236 (G4628gat, G4588gat);
nand NAND2_1237 (G4629gat, G4569gat, G4506gat);
not NOT1_1238 (G4630gat, G4569gat);
not NOT1_1239 (G4635gat, G4576gat);
nand NAND2_1240 (G4636gat, G4576gat, G4291gat);
not NOT1_1241 (G4640gat, G4581gat);
nand NAND2_1242 (G4641gat, G4581gat, G4461gat);
not NOT1_1243 (G4642gat, G4584gat);
nand NAND2_1244 (G4643gat, G4584gat, G4462gat);
nor NOR2_1245 (G4644gat, G4608gat, G4563gat);
and AND2_1246 (G4647gat, G4559gat, G2128gat);
and AND2_1247 (G4650gat, G4559gat, G2743gat);
and AND2_1248 (G4667gat, G4587gat, G4628gat);
nand NAND2_1249 (G4668gat, G4413gat, G4630gat);
not NOT1_1250 (G4669gat, G4616gat);
nand NAND2_1251 (G4670gat, G4616gat, G4239gat);
not NOT1_1252 (G4673gat, G4619gat);
nand NAND2_1253 (G4674gat, G4619gat, G4507gat);
nand NAND2_1254 (G4675gat, G4186gat, G4635gat);
not NOT1_1255 (G4676gat, G4623gat);
nand NAND2_1256 (G4677gat, G4623gat, G4558gat);
nand NAND2_1257 (G4678gat, G4365gat, G4640gat);
nand NAND2_1258 (G4679gat, G4368gat, G4642gat);
not NOT1_1259 (G4687gat, G4613gat);
nand NAND2_1260 (G4688gat, G4613gat, G4568gat);
nand NAND2_1261 (G4704gat, G4629gat, G4668gat);
nand NAND2_1262 (G4705gat, G4139gat, G4669gat);
not NOT1_1263 (G4706gat, G4656gat);
not NOT1_1264 (G4707gat, G4659gat);
nand NAND2_1265 (G4708gat, G4435gat, G4673gat);
nand NAND2_1266 (G4711gat, G4675gat, G4636gat);
nand NAND2_1267 (G4716gat, G4493gat, G4676gat);
nand NAND2_1268 (G4717gat, G4678gat, G4641gat);
nand NAND2_1269 (G4721gat, G4679gat, G4643gat);
not NOT1_1270 (G4726gat, G4664gat);
or OR3_1271 (G4727gat, G4647gat, G4650gat, G4350gat);
nor NOR3_1272 (G4730gat, G4647gat, G4650gat, G4350gat);
nand NAND2_1273 (G4733gat, G4479gat, G4687gat);
nand NAND2_1274 (G4740gat, G4705gat, G4670gat);
nand NAND2_1275 (G4743gat, G4708gat, G4674gat);
not NOT1_1276 (G4747gat, G4691gat);
nand NAND2_1277 (G4748gat, G4691gat, G4596gat);
not NOT1_1278 (G4749gat, G4694gat);
nand NAND2_1279 (G4750gat, G4694gat, G4597gat);
not NOT1_1280 (G4753gat, G4697gat);
nand NAND2_1281 (G4754gat, G4697gat, G4602gat);
not NOT1_1282 (G4755gat, G4700gat);
nand NAND2_1283 (G4756gat, G4700gat, G4603gat);
nand NAND2_1284 (G4757gat, G4716gat, G4677gat);
nand NAND2_1285 (G4769gat, G4733gat, G4688gat);
and AND2_1286 (G4772gat, G330gat, G4704gat);
not NOT1_1287 (G4775gat, G4721gat);
not NOT1_1288 (G4778gat, G4730gat);
nand NAND2_1289 (G4786gat, G4531gat, G4747gat);
nand NAND2_1290 (G4787gat, G4534gat, G4749gat);
nand NAND2_1291 (G4788gat, G4537gat, G4753gat);
nand NAND2_1292 (G4789gat, G4540gat, G4755gat);
and AND2_1293 (G4794gat, G4711gat, G2124gat);
and AND2_1294 (G4797gat, G4711gat, G2735gat);
and AND2_1295 (G4800gat, G4717gat, G2127gat);
and AND2_1296 (G4808gat, G4717gat, G4468gat);
and AND2_1297 (G4815gat, G4727gat, G4778gat);
not NOT1_1298 (G4816gat, G4769gat);
not NOT1_1299 (G4817gat, G4772gat);
nand NAND2_1300 (G4818gat, G4786gat, G4748gat);
nand NAND2_1301 (G4822gat, G4787gat, G4750gat);
nand NAND2_1302 (G4823gat, G4788gat, G4754gat);
nand NAND2_1303 (G4826gat, G4789gat, G4756gat);
nand NAND2_1304 (G4829gat, G4775gat, G4726gat);
not NOT1_1305 (G4830gat, G4775gat);
and AND2_1306 (G4831gat, G4743gat, G2122gat);
and AND2_1307 (G4838gat, G4757gat, G2126gat);
nand NAND2_1308 (G4859gat, G4772gat, G4816gat);
nand NAND2_1309 (G4860gat, G4769gat, G4817gat);
not NOT1_1310 (G4868gat, G4826gat);
not NOT1_1311 (G4870gat, G4805gat);
not NOT1_1312 (G4872gat, G4808gat);
nand NAND2_1313 (G4873gat, G4664gat, G4830gat);
or OR3_1314 (G4876gat, G4794gat, G4797gat, G4341gat);
nor NOR3_1315 (G4880gat, G4794gat, G4797gat, G4341gat);
not NOT1_1316 (G4885gat, G4812gat);
not NOT1_1317 (G4889gat, G4822gat);
nand NAND2_1318 (G4895gat, G4859gat, G4860gat);
not NOT1_1319 (G4896gat, G4844gat);
nand NAND2_1320 (G4897gat, G4844gat, G4706gat);
not NOT1_1321 (G4898gat, G4847gat);
nand NAND2_1322 (G4899gat, G4847gat, G4707gat);
nor NOR2_1323 (G4900gat, G4868gat, G4564gat);
and AND4_1324 (G4901gat, G4717gat, G4757gat, G4823gat, G4564gat);
not NOT1_1325 (G4902gat, G4850gat);
not NOT1_1326 (G4904gat, G4854gat);
nand NAND2_1327 (G4905gat, G4854gat, G4872gat);
nand NAND2_1328 (G4906gat, G4873gat, G4829gat);
and AND2_1329 (G4907gat, G4818gat, G2123gat);
and AND2_1330 (G4913gat, G4823gat, G2125gat);
and AND2_1331 (G4916gat, G4818gat, G4644gat);
not NOT1_1332 (G4920gat, G4880gat);
and AND2_1333 (G4921gat, G4895gat, G2184gat);
nand NAND2_1334 (G4924gat, G4656gat, G4896gat);
nand NAND2_1335 (G4925gat, G4659gat, G4898gat);
or OR2_1336 (G4926gat, G4900gat, G4901gat);
nand NAND2_1337 (G4928gat, G4889gat, G4870gat);
not NOT1_1338 (G4929gat, G4889gat);
nand NAND2_1339 (G4930gat, G4808gat, G4904gat);
not NOT1_1340 (G4931gat, G4906gat);
and AND2_1341 (G4944gat, G4876gat, G4920gat);
nand NAND2_1342 (G4946gat, G4924gat, G4897gat);
nand NAND2_1343 (G4949gat, G4925gat, G4899gat);
nand NAND2_1344 (G4950gat, G4916gat, G4902gat);
not NOT1_1345 (G4951gat, G4916gat);
nand NAND2_1346 (G4952gat, G4805gat, G4929gat);
nand NAND2_1347 (G4953gat, G4930gat, G4905gat);
and AND2_1348 (G4954gat, G4926gat, G2737gat);
and AND2_1349 (G4957gat, G4931gat, G2741gat);
or OR3_1350 (G4964gat, G2764gat, G2483gat, G4921gat);
nor NOR3_1351 (G4965gat, G2764gat, G2483gat, G4921gat);
not NOT1_1352 (G4968gat, G4949gat);
nand NAND2_1353 (G4969gat, G4850gat, G4951gat);
nand NAND2_1354 (G4970gat, G4952gat, G4928gat);
and AND2_1355 (G4973gat, G4953gat, G2739gat);
not NOT1_1356 (G4978gat, G4937gat);
not NOT1_1357 (G4979gat, G4940gat);
not NOT1_1358 (G4980gat, G4965gat);
nor NOR2_1359 (G4981gat, G4968gat, G4722gat);
and AND4_1360 (G4982gat, G4818gat, G4743gat, G4946gat, G4722gat);
nand NAND2_1361 (G4983gat, G4950gat, G4969gat);
not NOT1_1362 (G4984gat, G4970gat);
and AND2_1363 (G4985gat, G4946gat, G2121gat);
or OR3_1364 (G4988gat, G4913gat, G4954gat, G4344gat);
nor NOR3_1365 (G4991gat, G4913gat, G4954gat, G4344gat);
or OR3_1366 (G4996gat, G4800gat, G4957gat, G4347gat);
nor NOR3_1367 (G4999gat, G4800gat, G4957gat, G4347gat);
and AND2_1368 (G5002gat, G4964gat, G4980gat);
or OR2_1369 (G5007gat, G4981gat, G4982gat);
and AND2_1370 (G5010gat, G4983gat, G2731gat);
and AND2_1371 (G5013gat, G4984gat, G2733gat);
or OR3_1372 (G5018gat, G4838gat, G4973gat, G4475gat);
nor NOR3_1373 (G5021gat, G4838gat, G4973gat, G4475gat);
not NOT1_1374 (G5026gat, G4991gat);
not NOT1_1375 (G5029gat, G4999gat);
and AND2_1376 (G5030gat, G5007gat, G2729gat);
and AND2_1377 (G5045gat, G4988gat, G5026gat);
not NOT1_1378 (G5046gat, G5021gat);
and AND2_1379 (G5047gat, G4996gat, G5029gat);
or OR3_1380 (G5050gat, G4831gat, G5010gat, G4472gat);
nor NOR3_1381 (G5055gat, G4831gat, G5010gat, G4472gat);
or OR3_1382 (G5058gat, G4907gat, G5013gat, G4338gat);
nor NOR3_1383 (G5061gat, G4907gat, G5013gat, G4338gat);
and AND4_1384 (G5066gat, G4730gat, G4999gat, G5021gat, G4991gat);
and AND2_1385 (G5078gat, G5018gat, G5046gat);
or OR3_1386 (G5080gat, G4985gat, G5030gat, G4335gat);
nor NOR3_1387 (G5085gat, G4985gat, G5030gat, G4335gat);
nand NAND2_1388 (G5094gat, G5039gat, G4885gat);
not NOT1_1389 (G5095gat, G5039gat);
not NOT1_1390 (G5097gat, G5042gat);
and AND2_1391 (G5102gat, G5050gat, G5050gat);
not NOT1_1392 (G5103gat, G5061gat);
nand NAND2_1393 (G5108gat, G4812gat, G5095gat);
not NOT1_1394 (G5109gat, G5070gat);
nand NAND2_1395 (G5110gat, G5070gat, G5097gat);
and AND2_1396 (G5114gat, G5050gat, G1461gat);
and AND2_1397 (G5120gat, G5080gat, G5080gat);
and AND2_1398 (G5121gat, G5058gat, G5103gat);
nand NAND2_1399 (G5122gat, G5094gat, G5108gat);
nand NAND2_1400 (G5125gat, G5042gat, G5109gat);
and AND2_1401 (G5128gat, G1461gat, G5080gat);
and AND4_1402 (G5133gat, G4880gat, G5061gat, G5055gat, G5085gat);
and AND3_1403 (G5136gat, G5055gat, G5085gat, G1464gat);
nand NAND2_1404 (G5145gat, G5125gat, G5110gat);
not NOT1_1405 (G5159gat, G5117gat);
and AND2_1406 (G5166gat, G5066gat, G5133gat);
and AND2_1407 (G5173gat, G5066gat, G5133gat);
not NOT1_1408 (G5182gat, G5139gat);
nand NAND2_1409 (G5183gat, G5139gat, G5159gat);
not NOT1_1410 (G5192gat, G5166gat);
nor NOR2_1411 (G5193gat, G5136gat, G5173gat);
nand NAND2_1412 (G5196gat, G5151gat, G4978gat);
not NOT1_1413 (G5197gat, G5151gat);
nand NAND2_1414 (G5198gat, G5154gat, G4979gat);
not NOT1_1415 (G5199gat, G5154gat);
not NOT1_1416 (G5201gat, G5160gat);
not NOT1_1417 (G5203gat, G5163gat);
nand NAND2_1418 (G5212gat, G5117gat, G5182gat);
and AND2_1419 (G5215gat, G213gat, G5193gat);
not NOT1_1420 (G5217gat, G5174gat);
not NOT1_1421 (G5219gat, G5177gat);
nand NAND2_1422 (G5220gat, G4937gat, G5197gat);
nand NAND2_1423 (G5221gat, G4940gat, G5199gat);
not NOT1_1424 (G5222gat, G5184gat);
nand NAND2_1425 (G5223gat, G5184gat, G5201gat);
nand NAND2_1426 (G5224gat, G5188gat, G5203gat);
not NOT1_1427 (G5225gat, G5188gat);
nand NAND2_1428 (G5228gat, G5183gat, G5212gat);
not NOT1_1429 (G5231gat, G5215gat);
nand NAND2_1430 (G5232gat, G5205gat, G5217gat);
not NOT1_1431 (G5233gat, G5205gat);
nand NAND2_1432 (G5234gat, G5209gat, G5219gat);
not NOT1_1433 (G5235gat, G5209gat);
nand NAND2_1434 (G5236gat, G5196gat, G5220gat);
nand NAND2_1435 (G5240gat, G5198gat, G5221gat);
nand NAND2_1436 (G5242gat, G5160gat, G5222gat);
nand NAND2_1437 (G5243gat, G5163gat, G5225gat);
nand NAND2_1438 (G5245gat, G5174gat, G5233gat);
nand NAND2_1439 (G5246gat, G5177gat, G5235gat);
not NOT1_1440 (G5250gat, G5240gat);
not NOT1_1441 (G5253gat, G5228gat);
nand NAND2_1442 (G5254gat, G5242gat, G5223gat);
nand NAND2_1443 (G5257gat, G5243gat, G5224gat);
nand NAND2_1444 (G5258gat, G5232gat, G5245gat);
nand NAND2_1445 (G5261gat, G5234gat, G5246gat);
not NOT1_1446 (G5266gat, G5257gat);
and AND3_1447 (G5277gat, G5236gat, G5254gat, G2307gat);
and AND3_1448 (G5278gat, G5250gat, G5254gat, G2310gat);
not NOT1_1449 (G5279gat, G5261gat);
not NOT1_1450 (G5283gat, G5269gat);
nand NAND2_1451 (G5284gat, G5269gat, G5253gat);
and AND3_1452 (G5285gat, G5236gat, G5266gat, G2310gat);
and AND3_1453 (G5286gat, G5250gat, G5266gat, G2307gat);
nand NAND2_1454 (G5295gat, G5228gat, G5283gat);
or OR4_1455 (G5298gat, G5277gat, G5285gat, G5278gat, G5286gat);
nand NAND2_1456 (G5309gat, G5295gat, G5284gat);
not NOT1_1457 (G5312gat, G5292gat);
not NOT1_1458 (G5313gat, G5289gat);
not NOT1_1459 (G5322gat, G5306gat);
not NOT1_1460 (G5323gat, G5303gat);
nand NAND2_1461 (G5340gat, G5324gat, G5323gat);
nand NAND2_1462 (G5341gat, G5327gat, G5322gat);
not NOT1_1463 (G5344gat, G5327gat);
not NOT1_1464 (G5345gat, G5324gat);
nand NAND2_1465 (G5348gat, G5332gat, G5313gat);
nand NAND2_1466 (G5349gat, G5335gat, G5312gat);
nand NAND2_1467 (G5350gat, G5303gat, G5345gat);
nand NAND2_1468 (G5351gat, G5306gat, G5344gat);
not NOT1_1469 (G5352gat, G5335gat);
not NOT1_1470 (G5353gat, G5332gat);
nand NAND2_1471 (G5354gat, G5289gat, G5353gat);
nand NAND2_1472 (G5355gat, G5292gat, G5352gat);
nand NAND2_1473 (G5356gat, G5350gat, G5340gat);
nand NAND2_1474 (G5357gat, G5351gat, G5341gat);
nand NAND2_1475 (G5358gat, G5348gat, G5354gat);
nand NAND2_1476 (G5359gat, G5349gat, G5355gat);
and AND2_1477 (G5360gat, G5356gat, G5357gat);
nand NAND2_1478 (G5361gat_enc, G5358gat, G5359gat);
xor XOR2_1479 (nXOR0, G1gat, keyinput0);
xor XOR2_1480 (nXOR1, G13gat, keyinput1);
xor XOR2_1481 (nXOR2, G20gat, keyinput2);
xor XOR2_1482 (nXOR3, G33gat, keyinput3);
xor XOR2_1483 (nXOR4, G41gat, keyinput4);
xor XOR2_1484 (nXOR5, G45gat, keyinput5);
xor XOR2_1485 (nXOR6, G50gat, keyinput6);
xor XOR2_1486 (nXOR7, G58gat, keyinput7);
not NOT1_1487 (not_keyinp0, keyinput0);
not NOT1_1488 (not_keyinp1, keyinput1);
not NOT1_1489 (not_keyinp2, keyinput2);
not NOT1_1490 (not_keyinp3, keyinput3);
not NOT1_1491 (not_keyinp4, keyinput4);
not NOT1_1492 (not_keyinp5, keyinput5);
not NOT1_1493 (not_keyinp6, keyinput6);
not NOT1_1494 (not_keyinp7, keyinput7);
nor NOR8_1495 (flipSig, nXOR0, nXOR1, nXOR2, nXOR3, nXOR4, nXOR5, nXOR6, nXOR7);
and AND8_1496 (maskSig, keyinput0, not_keyinp1, keyinput2, keyinput3, not_keyinp4, not_keyinp5, keyinput6, not_keyinp7);
not NOT1_1497 (not_mask, maskSig);
and AND2_1498 (flip_mask, flipSig, not_mask);
xor XOR2_1499 (G5361gat, flip_mask, G5361gat_enc);

endmodule