module ttlock(keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,n6123);

input keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31;
output n6123;
wire n_0,wire1316,wire1318,wire1419,wire1420,wire1328,wire1499,wire1500,wire1320,wire1322,wire1503,wire1504,wire1300,wire1302,wire1381,wire1385,wire1357,wire1393,wire1332,wire1365,wire1361,wire1415,wire1416,wire1308,wire1310,wire1373,wire1375,wire1405,wire1407,wire1312,wire1314,wire1389,wire1391,wire1508,wire1509,wire1340,wire1342,wire1324,wire1326,wire1304,wire1306,wire1423,wire1424,wire1401,wire1403,wire1369,wire1371,wire1397,wire1399,wire1377,wire1379,wire1336,wire1338,wire1353,wire1355,wire1285,wire1286,wire1317,wire1421,wire1329,wire1330,wire1501,wire1321,wire1505,wire1301,wire1382,wire1383,wire1386,wire1387,wire1358,wire1359,wire1394,wire1395,wire1333,wire1334,wire1366,wire1367,wire1362,wire1363,wire1417,wire1309,wire1374,wire1406,wire1313,wire1390,wire1510,wire1341,wire1325,wire1305,wire1425,wire1402,wire1370,wire1398,wire1378,wire1337,wire1354,wire1287,wire1319,wire1422,wire1331,wire1502,wire1323,wire1506,wire1303,wire1384,wire1388,wire1360,wire1396,wire1335,wire1368,wire1364,wire1418,wire1311,wire1376,wire1408,wire1315,wire1392,wire1511,wire1343,wire1327,wire1307,wire1426,wire1404,wire1372,wire1400,wire1380,wire1339,wire1356,n_73,n_31,n_69,n_5,n_72,n_4,n_78,n_48,n_47,n_54,n_45,n_68,n_52,n_53,n_32,n_76,n_50,n_42,n_75,n_46,n_1,n_66,n_71,n_77,n_30,n_43,n_51,n_44,n_49,n_67,n_56,wire1288,wire1284,wire1290,wire1280,wire1282,wire1283,wire1281,wire1289,n_98,n_99,n_95,n_104,n_101,n_100,n_103,n_96,wire1246,wire1245,n_122,n_123,wire1222,n_1429,wire66,wire67,wire68,wire69;

not NOT1_1 (n_0, keyinput0);
not NOT1_2 (wire1316, keyinput1);
and AND2_3 (wire1318, keyinput1, n290);
or OR2_4 (wire1419, n239, keyinput2);
and AND2_5 (wire1420, n239, keyinput2);
not NOT1_6 (wire1328, keyinput3);
and AND2_7 (wire1499, n222, keyinput4);
or OR2_8 (wire1500, n222, keyinput4);
not NOT1_9 (wire1320, keyinput5);
and AND2_10 (wire1322, keyinput5, n273);
and AND2_11 (wire1503, n205, keyinput6);
or OR2_12 (wire1504, n205, keyinput6);
not NOT1_13 (wire1300, keyinput7);
and AND2_14 (wire1302, keyinput7, n324);
not NOT1_15 (wire1381, keyinput8);
not NOT1_16 (wire1385, keyinput9);
not NOT1_17 (wire1357, keyinput10);
not NOT1_18 (wire1393, keyinput11);
not NOT1_19 (wire1332, keyinput12);
not NOT1_20 (wire1365, keyinput13);
not NOT1_21 (wire1361, keyinput14);
or OR2_22 (wire1415, n392, keyinput15);
and AND2_23 (wire1416, n392, keyinput15);
not NOT1_24 (wire1308, keyinput16);
and AND2_25 (wire1310, keyinput16, n120);
not NOT1_26 (wire1373, keyinput17);
and AND2_27 (wire1375, keyinput17, n409);
not NOT1_28 (wire1405, keyinput18);
and AND2_29 (wire1407, keyinput18, n103);
not NOT1_30 (wire1312, keyinput19);
and AND2_31 (wire1314, keyinput19, n426);
not NOT1_32 (wire1389, keyinput20);
and AND2_33 (wire1391, keyinput20, n86);
and AND2_34 (wire1508, n443, keyinput21);
or OR2_35 (wire1509, n443, keyinput21);
not NOT1_36 (wire1340, keyinput22);
and AND2_37 (wire1342, keyinput22, n69);
not NOT1_38 (wire1324, keyinput23);
and AND2_39 (wire1326, keyinput23, n460);
not NOT1_40 (wire1304, keyinput24);
and AND2_41 (wire1306, keyinput24, n52);
and AND2_42 (wire1423, n477, keyinput25);
or OR2_43 (wire1424, n477, keyinput25);
not NOT1_44 (wire1401, keyinput26);
and AND2_45 (wire1403, keyinput26, n35);
not NOT1_46 (wire1369, keyinput27);
and AND2_47 (wire1371, keyinput27, n494);
not NOT1_48 (wire1397, keyinput28);
and AND2_49 (wire1399, keyinput28, n18);
not NOT1_50 (wire1377, keyinput29);
and AND2_51 (wire1379, keyinput29, n511);
not NOT1_52 (wire1336, keyinput30);
and AND2_53 (wire1338, keyinput30, n528);
not NOT1_54 (wire1353, keyinput31);
and AND2_55 (wire1355, keyinput31, n1);
and AND2_56 (wire1285, n_0, n256);
and AND2_57 (wire1286, n_97, keyinput0);
and AND2_58 (wire1317, wire1316, n_155);
not NOT1_59 (wire1421, wire1420);
and AND2_60 (wire1329, wire1328, n307);
and AND2_61 (wire1330, keyinput3, n_207);
not NOT1_62 (wire1501, wire1500);
and AND2_63 (wire1321, wire1320, n_2);
not NOT1_64 (wire1505, wire1504);
and AND2_65 (wire1301, wire1300, n_22);
and AND2_66 (wire1382, wire1381, n188);
and AND2_67 (wire1383, keyinput8, n_25);
and AND2_68 (wire1386, wire1385, n341);
and AND2_69 (wire1387, keyinput9, n_21);
and AND2_70 (wire1358, wire1357, n171);
and AND2_71 (wire1359, keyinput10, n_9);
and AND2_72 (wire1394, wire1393, n358);
and AND2_73 (wire1395, keyinput11, n_14);
and AND2_74 (wire1333, wire1332, n154);
and AND2_75 (wire1334, keyinput12, n_20);
and AND2_76 (wire1366, wire1365, n375);
and AND2_77 (wire1367, keyinput13, n_27);
and AND2_78 (wire1362, wire1361, n137);
and AND2_79 (wire1363, keyinput14, n_6);
not NOT1_80 (wire1417, wire1416);
and AND2_81 (wire1309, wire1308, n_11);
and AND2_82 (wire1374, wire1373, n_16);
and AND2_83 (wire1406, wire1405, n_41);
and AND2_84 (wire1313, wire1312, n_74);
and AND2_85 (wire1390, wire1389, n_24);
not NOT1_86 (wire1510, wire1509);
and AND2_87 (wire1341, wire1340, n_29);
and AND2_88 (wire1325, wire1324, n_70);
and AND2_89 (wire1305, wire1304, n_13);
not NOT1_90 (wire1425, wire1424);
and AND2_91 (wire1402, wire1401, n_26);
and AND2_92 (wire1370, wire1369, n_10);
and AND2_93 (wire1398, wire1397, n_18);
and AND2_94 (wire1378, wire1377, n_17);
and AND2_95 (wire1337, wire1336, n_7);
and AND2_96 (wire1354, wire1353, n_55);
or OR2_97 (wire1287, wire1286, wire1285);
or OR2_98 (wire1319, wire1318, wire1317);
and AND2_99 (wire1422, wire1421, wire1419);
or OR2_100 (wire1331, wire1330, wire1329);
or OR2_101 (wire1502, wire1501, wire1499);
or OR2_102 (wire1323, wire1322, wire1321);
or OR2_103 (wire1506, wire1505, wire1503);
or OR2_104 (wire1303, wire1302, wire1301);
or OR2_105 (wire1384, wire1383, wire1382);
or OR2_106 (wire1388, wire1387, wire1386);
or OR2_107 (wire1360, wire1359, wire1358);
or OR2_108 (wire1396, wire1395, wire1394);
or OR2_109 (wire1335, wire1334, wire1333);
or OR2_110 (wire1368, wire1367, wire1366);
or OR2_111 (wire1364, wire1363, wire1362);
and AND2_112 (wire1418, wire1417, wire1415);
or OR2_113 (wire1311, wire1310, wire1309);
or OR2_114 (wire1376, wire1375, wire1374);
or OR2_115 (wire1408, wire1407, wire1406);
or OR2_116 (wire1315, wire1314, wire1313);
or OR2_117 (wire1392, wire1391, wire1390);
or OR2_118 (wire1511, wire1510, wire1508);
or OR2_119 (wire1343, wire1342, wire1341);
or OR2_120 (wire1327, wire1326, wire1325);
or OR2_121 (wire1307, wire1306, wire1305);
or OR2_122 (wire1426, wire1425, wire1423);
or OR2_123 (wire1404, wire1403, wire1402);
or OR2_124 (wire1372, wire1371, wire1370);
or OR2_125 (wire1400, wire1399, wire1398);
or OR2_126 (wire1380, wire1379, wire1378);
or OR2_127 (wire1339, wire1338, wire1337);
or OR2_128 (wire1356, wire1355, wire1354);
not NOT1_129 (n_73, wire1319);
not NOT1_130 (n_31, wire1422);
not NOT1_131 (n_69, wire1331);
not NOT1_132 (n_5, wire1502);
not NOT1_133 (n_72, wire1323);
not NOT1_134 (n_4, wire1506);
not NOT1_135 (n_78, wire1303);
not NOT1_136 (n_48, wire1384);
not NOT1_137 (n_47, wire1388);
not NOT1_138 (n_54, wire1360);
not NOT1_139 (n_45, wire1396);
not NOT1_140 (n_68, wire1335);
not NOT1_141 (n_52, wire1368);
not NOT1_142 (n_53, wire1364);
not NOT1_143 (n_32, wire1418);
not NOT1_144 (n_76, wire1311);
not NOT1_145 (n_50, wire1376);
not NOT1_146 (n_42, wire1408);
not NOT1_147 (n_75, wire1315);
not NOT1_148 (n_46, wire1392);
not NOT1_149 (n_1, wire1511);
not NOT1_150 (n_66, wire1343);
not NOT1_151 (n_71, wire1327);
not NOT1_152 (n_77, wire1307);
not NOT1_153 (n_30, wire1426);
not NOT1_154 (n_43, wire1404);
not NOT1_155 (n_51, wire1372);
not NOT1_156 (n_44, wire1400);
not NOT1_157 (n_49, wire1380);
not NOT1_158 (n_67, wire1339);
not NOT1_159 (n_56, wire1356);
or OR2_160 (wire1288, wire1287, n_73);
or OR4_161 (wire1284, n_72, n_78, n_4, n_5);
and AND4_162 (wire1290, n_48, n_54, n_45, n_47);
and AND4_163 (wire1280, n_53, n_68, n_52, n_32);
or OR4_164 (wire1282, n_75, n_42, n_50, n_76);
or OR4_165 (wire1283, n_66, n_46, n_71, n_1);
or OR4_166 (wire1281, n_51, n_77, n_43, n_30);
or OR4_167 (wire1289, n_56, n_67, n_49, n_44);
not NOT1_168 (n_98, wire1288);
not NOT1_169 (n_99, wire1284);
not NOT1_170 (n_95, wire1290);
not NOT1_171 (n_104, wire1280);
not NOT1_172 (n_101, wire1282);
not NOT1_173 (n_100, wire1283);
not NOT1_174 (n_103, wire1281);
not NOT1_175 (n_96, wire1289);
and AND4_176 (wire1246, n_99, n_98, n_69, n_31);
and AND4_177 (wire1245, n_101, n_96, n_100, n_103);
not NOT1_178 (n_122, wire1246);
not NOT1_179 (n_123, wire1245);
or OR4_180 (wire1222, n_123, n_122, n_95, n_104);
not NOT1_181 (n_1429, wire1222);
or OR2_182 (wire66, n_1430, n_1429);
and AND2_183 (wire67, n_1430, n_1429);
not NOT1_184 (wire68, wire67);
and AND2_185 (wire69, wire68, wire66);
not NOT1_186 (n6123, wire69);

endmodule