module DFF(Q, clk, D);
input D;
input clk;
output Q;
always @(clk)
begin
  Q <= D;
end
endmodule


module c1355_libar_32k(G1gat,G8gat,G15gat,G22gat,G29gat,G36gat,G43gat,G50gat,G57gat,G64gat,G71gat,G78gat,G85gat,G92gat,G99gat,G106gat,G113gat,G120gat,G127gat,G134gat,G141gat,G148gat,G155gat,G162gat,G169gat,G176gat,G183gat,G190gat,G197gat,G204gat,G211gat,G218gat,G225gat,G226gat,G227gat,G228gat,G229gat,G230gat,G231gat,G232gat,G233gat,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,G1324gat,G1325gat,G1326gat,G1327gat,G1328gat,G1329gat,G1330gat,G1331gat,G1332gat,G1333gat,G1334gat,G1335gat,G1336gat,G1337gat,G1338gat,G1339gat,G1340gat,G1341gat,G1342gat,G1343gat,G1344gat,G1345gat,G1346gat,G1347gat,G1348gat,G1349gat,G1350gat,G1351gat,G1352gat,G1353gat,G1354gat,G1355gat);

input G1gat,G8gat,G15gat,G22gat,G29gat,G36gat,G43gat,G50gat,G57gat,G64gat,G71gat,G78gat,G85gat,G92gat,G99gat,G106gat,G113gat,G120gat,G127gat,G134gat,G141gat,G148gat,G155gat,G162gat,G169gat,G176gat,G183gat,G190gat,G197gat,G204gat,G211gat,G218gat,G225gat,G226gat,G227gat,G228gat,G229gat,G230gat,G231gat,G232gat,G233gat,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31;
output G1324gat,G1325gat,G1326gat,G1327gat,G1328gat,G1329gat,G1330gat,G1331gat,G1332gat,G1333gat,G1334gat,G1335gat,G1336gat,G1337gat,G1338gat,G1339gat,G1340gat,G1341gat,G1342gat,G1343gat,G1344gat,G1345gat,G1346gat,G1347gat,G1348gat,G1349gat,G1350gat,G1351gat,G1352gat,G1353gat,G1354gat,G1355gat;
wire G242gat,G245gat,G248gat_enc,CLK11,LIBAR11,G248gat,G251gat_enc,G251gat,G254gat_enc,CLK10,LIBAR10,G254gat,G257gat,G260gat_enc,G260gat,G263gat,G266gat,G269gat,G272gat,G275gat_enc,CLK9,LIBAR9,G275gat,G278gat_enc,G278gat,G281gat_enc,CLK8,LIBAR8,G281gat,G284gat_enc,G284gat,G287gat_enc,CLK7,LIBAR7,G287gat,G290gat_enc,CLK6,LIBAR6,G290gat,G293gat_enc,G293gat,G296gat,G299gat_enc,CLK5,LIBAR5,G299gat,G302gat,G305gat_enc,CLK4,LIBAR4,G305gat,G308gat_enc,CLK3,LIBAR3,G308gat,G311gat_enc,CLK2,LIBAR2,G311gat,G314gat_enc,G314gat,G317gat,G320gat,G323gat,G326gat_enc,CLK1,LIBAR1,G326gat,G329gat_enc,G329gat,G332gat,G335gat_enc,G335gat,G338gat_enc,G338gat,G341gat_enc,G341gat,G344gat,G347gat_enc,G347gat,G350gat,G353gat_enc,G353gat,G356gat,G359gat_enc,G359gat,G362gat_enc,G362gat,G363gat,G364gat,G365gat,G366gat_enc,G366gat,G367gat_enc,G367gat,G368gat_enc,G368gat,G369gat_enc,G369gat,G370gat_enc,G370gat,G371gat_enc,G371gat,G372gat,G373gat,G374gat_enc,G374gat,G375gat,G376gat,G377gat,G378gat,G379gat,G380gat,G381gat,G382gat,G383gat,G384gat,G385gat,G386gat,G387gat,G388gat,G389gat,G390gat,G391gat,G392gat,G393gat,G394gat,G395gat,G396gat,G397gat,G398gat,G399gat,G400gat,G401gat,G402gat,G403gat,G404gat,G405gat,G406gat,G407gat,G408gat,G409gat,G410gat,G411gat,G412gat,G413gat,G414gat,G415gat,G416gat,G417gat,G418gat,G419gat,G420gat,G421gat,G422gat,G423gat,G424gat,G425gat,G426gat,G429gat,G432gat,G435gat,G438gat,G441gat,G444gat,G447gat,G450gat,G453gat,G456gat,G459gat,G462gat,G465gat,G468gat,G471gat,G474gat,G477gat,G480gat,G483gat,G486gat,G489gat,G492gat,G495gat,G498gat,G501gat,G504gat,G507gat,G510gat,G513gat,G516gat,G519gat,G522gat,G525gat,G528gat,G531gat,G534gat,G537gat,G540gat,G543gat,G546gat,G549gat,G552gat,G555gat,G558gat,G561gat,G564gat,G567gat,G570gat,G571gat,G572gat,G573gat,G574gat,G575gat,G576gat,G577gat,G578gat,G579gat,G580gat,G581gat,G582gat,G583gat,G584gat,G585gat,G586gat,G587gat,G588gat,G589gat,G590gat,G591gat,G592gat,G593gat,G594gat,G595gat,G596gat,G597gat,G598gat,G599gat,G600gat,G601gat,G602gat,G607gat,G612gat,G617gat,G622gat,G627gat,G632gat,G637gat,G642gat,G645gat,G648gat,G651gat,G654gat,G657gat,G660gat,G663gat,G666gat,G669gat,G672gat,G675gat,G678gat,G681gat,G684gat,G687gat,G690gat,G691gat,G692gat,G693gat,G694gat,G695gat,G696gat,G697gat,G698gat,G699gat,G700gat,G701gat,G702gat,G703gat,G704gat,G705gat,G706gat,G709gat,G712gat,G715gat,G718gat,G721gat,G724gat,G727gat,G730gat,G733gat,G736gat,G739gat,G742gat,G745gat,G748gat,G751gat,G754gat,G755gat,G756gat,G757gat,G758gat,G759gat,G760gat,G761gat,G762gat,G763gat,G764gat,G765gat,G766gat,G767gat,G768gat,G769gat,G770gat,G773gat,G776gat,G779gat,G782gat,G785gat,G788gat,G791gat,G794gat,G797gat,G800gat,G803gat,G806gat,G809gat,G812gat,G815gat,G818gat,G819gat,G820gat,G821gat,G822gat,G823gat,G824gat,G825gat,G826gat,G827gat,G828gat,G829gat,G830gat,G831gat,G832gat,G833gat,G834gat,G847gat,G860gat,G873gat,G886gat,G899gat,G912gat,G925gat,G938gat,G939gat,G940gat,G941gat,G942gat,G943gat,G944gat,G945gat,G946gat,G947gat,G948gat,G949gat,G950gat,G951gat,G952gat,G953gat,G954gat,G955gat,G956gat,G957gat,G958gat,G959gat,G960gat,G961gat,G962gat,G963gat,G964gat,G965gat,G966gat,G967gat,G968gat,G969gat,G970gat,G971gat,G972gat,G973gat,G974gat,G975gat,G976gat,G977gat,G978gat,G979gat,G980gat,G981gat,G982gat,G983gat,G984gat,G985gat,G986gat,G991gat,G996gat,G1001gat,G1006gat,G1011gat,G1016gat,G1021gat,G1026gat,G1031gat,G1036gat,G1039gat,G1042gat,G1045gat,G1048gat,G1051gat,G1054gat,G1057gat,G1060gat,G1063gat,G1066gat,G1069gat,G1072gat,G1075gat,G1078gat,G1081gat,G1084gat,G1087gat,G1090gat,G1093gat,G1096gat,G1099gat,G1102gat,G1105gat,G1108gat,G1111gat,G1114gat,G1117gat,G1120gat,G1123gat,G1126gat,G1129gat,G1132gat,G1135gat,G1138gat,G1141gat,G1144gat,G1147gat,G1150gat,G1153gat,G1156gat,G1159gat,G1162gat,G1165gat,G1168gat,G1171gat,G1174gat,G1177gat,G1180gat,G1183gat,G1186gat,G1189gat,G1192gat,G1195gat,G1198gat,G1201gat,G1204gat,G1207gat,G1210gat,G1213gat,G1216gat,G1219gat,G1222gat,G1225gat,G1228gat,G1229gat,G1230gat,G1231gat,G1232gat,G1233gat,G1234gat,G1235gat,G1236gat,G1237gat,G1238gat,G1239gat,G1240gat,G1241gat,G1242gat,G1243gat,G1244gat,G1245gat,G1246gat,G1247gat,G1248gat,G1249gat,G1250gat,G1251gat,G1252gat,G1253gat,G1254gat,G1255gat,G1256gat,G1257gat,G1258gat,G1259gat,G1260gat,G1261gat,G1262gat,G1263gat,G1264gat,G1265gat,G1266gat,G1267gat,G1268gat,G1269gat,G1270gat,G1271gat,G1272gat,G1273gat,G1274gat,G1275gat,G1276gat,G1277gat,G1278gat,G1279gat,G1280gat,G1281gat,G1282gat,G1283gat,G1284gat,G1285gat,G1286gat,G1287gat,G1288gat,G1289gat,G1290gat,G1291gat,G1292gat,G1293gat,G1294gat,G1295gat,G1296gat,G1297gat,G1298gat,G1299gat,G1300gat,G1301gat,G1302gat,G1303gat,G1304gat,G1305gat,G1306gat,G1307gat,G1308gat,G1309gat,G1310gat,G1311gat,G1312gat,G1313gat,G1314gat,G1315gat,G1316gat,G1317gat,G1318gat,G1319gat,G1320gat,G1321gat,G1322gat,G1323gat;

and AND2_1 (G242gat, G225gat, G233gat);
and AND2_2 (G245gat, G226gat, G233gat);
and AND2_3 (G248gat_enc, G227gat, G233gat);
nor NOR2_4 (CLK11, G248gat_enc, G245gat);
dff DFF2_5 (LIBAR11, CLK11, keyinput0);
xnor XNOR2_6 (G248gat, LIBAR11, G248gat_enc);
and AND2_7 (G251gat_enc, G228gat, G233gat);
xor XOR2_8 (G251gat, keyinput1, G251gat_enc);
and AND2_9 (G254gat_enc, G229gat, G233gat);
nor NOR2_10 (CLK10, G254gat_enc, G251gat);
dff DFF2_11 (LIBAR10, CLK10, keyinput2);
xor XOR2_12 (G254gat, LIBAR10, G254gat_enc);
and AND2_13 (G257gat, G230gat, G233gat);
and AND2_14 (G260gat_enc, G231gat, G233gat);
xnor XNOR2_15 (G260gat, keyinput3, G260gat_enc);
and AND2_16 (G263gat, G232gat, G233gat);
nand NAND2_17 (G266gat, G1gat, G8gat);
nand NAND2_18 (G269gat, G15gat, G22gat);
nand NAND2_19 (G272gat, G29gat, G36gat);
nand NAND2_20 (G275gat_enc, G43gat, G50gat);
nor NOR2_21 (CLK9, G275gat_enc, G272gat);
dff DFF2_22 (LIBAR9, CLK9, keyinput4);
xnor XNOR2_23 (G275gat, LIBAR9, G275gat_enc);
nand NAND2_24 (G278gat_enc, G57gat, G64gat);
xor XOR2_25 (G278gat, keyinput5, G278gat_enc);
nand NAND2_26 (G281gat_enc, G71gat, G78gat);
nor NOR2_27 (CLK8, G281gat_enc, G278gat);
dff DFF2_28 (LIBAR8, CLK8, keyinput6);
xor XOR2_29 (G281gat, LIBAR8, G281gat_enc);
nand NAND2_30 (G284gat_enc, G85gat, G92gat);
xor XOR2_31 (G284gat, keyinput7, G284gat_enc);
nand NAND2_32 (G287gat_enc, G99gat, G106gat);
nor NOR2_33 (CLK7, G287gat_enc, G284gat);
dff DFF2_34 (LIBAR7, CLK7, keyinput8);
xnor XNOR2_35 (G287gat, LIBAR7, G287gat_enc);
nand NAND2_36 (G290gat_enc, G113gat, G120gat);
nor NOR2_37 (CLK6, G290gat_enc, G287gat);
dff DFF2_38 (LIBAR6, CLK6, keyinput9);
xnor XNOR2_39 (G290gat, LIBAR6, G290gat_enc);
nand NAND2_40 (G293gat_enc, G127gat, G134gat);
xnor XNOR2_41 (G293gat, keyinput10, G293gat_enc);
nand NAND2_42 (G296gat, G141gat, G148gat);
nand NAND2_43 (G299gat_enc, G155gat, G162gat);
nor NOR2_44 (CLK5, G299gat_enc, G296gat);
dff DFF2_45 (LIBAR5, CLK5, keyinput11);
xnor XNOR2_46 (G299gat, LIBAR5, G299gat_enc);
nand NAND2_47 (G302gat, G169gat, G176gat);
nand NAND2_48 (G305gat_enc, G183gat, G190gat);
nor NOR2_49 (CLK4, G305gat_enc, G302gat);
dff DFF2_50 (LIBAR4, CLK4, keyinput12);
xnor XNOR2_51 (G305gat, LIBAR4, G305gat_enc);
nand NAND2_52 (G308gat_enc, G197gat, G204gat);
nor NOR2_53 (CLK3, G308gat_enc, G305gat);
dff DFF2_54 (LIBAR3, CLK3, keyinput13);
xor XOR2_55 (G308gat, LIBAR3, G308gat_enc);
nand NAND2_56 (G311gat_enc, G211gat, G218gat);
nor NOR2_57 (CLK2, G311gat_enc, G308gat);
dff DFF2_58 (LIBAR2, CLK2, keyinput14);
xnor XNOR2_59 (G311gat, LIBAR2, G311gat_enc);
nand NAND2_60 (G314gat_enc, G1gat, G29gat);
xor XOR2_61 (G314gat, keyinput15, G314gat_enc);
nand NAND2_62 (G317gat, G57gat, G85gat);
nand NAND2_63 (G320gat, G8gat, G36gat);
nand NAND2_64 (G323gat, G64gat, G92gat);
nand NAND2_65 (G326gat_enc, G15gat, G43gat);
nor NOR2_66 (CLK1, G326gat_enc, G323gat);
dff DFF2_67 (LIBAR1, CLK1, keyinput16);
xnor XNOR2_68 (G326gat, LIBAR1, G326gat_enc);
nand NAND2_69 (G329gat_enc, G71gat, G99gat);
xor XOR2_70 (G329gat, keyinput17, G329gat_enc);
nand NAND2_71 (G332gat, G22gat, G50gat);
nand NAND2_72 (G335gat_enc, G78gat, G106gat);
xnor XNOR2_73 (G335gat, keyinput18, G335gat_enc);
nand NAND2_74 (G338gat_enc, G113gat, G141gat);
xor XOR2_75 (G338gat, keyinput19, G338gat_enc);
nand NAND2_76 (G341gat_enc, G169gat, G197gat);
xnor XNOR2_77 (G341gat, keyinput20, G341gat_enc);
nand NAND2_78 (G344gat, G120gat, G148gat);
nand NAND2_79 (G347gat_enc, G176gat, G204gat);
xnor XNOR2_80 (G347gat, keyinput21, G347gat_enc);
nand NAND2_81 (G350gat, G127gat, G155gat);
nand NAND2_82 (G353gat_enc, G183gat, G211gat);
xnor XNOR2_83 (G353gat, keyinput22, G353gat_enc);
nand NAND2_84 (G356gat, G134gat, G162gat);
nand NAND2_85 (G359gat_enc, G190gat, G218gat);
xnor XNOR2_86 (G359gat, keyinput23, G359gat_enc);
nand NAND2_87 (G362gat_enc, G1gat, G266gat);
xor XOR2_88 (G362gat, keyinput24, G362gat_enc);
nand NAND2_89 (G363gat, G8gat, G266gat);
nand NAND2_90 (G364gat, G15gat, G269gat);
nand NAND2_91 (G365gat, G22gat, G269gat);
nand NAND2_92 (G366gat_enc, G29gat, G272gat);
xnor XNOR2_93 (G366gat, keyinput25, G366gat_enc);
nand NAND2_94 (G367gat_enc, G36gat, G272gat);
xor XOR2_95 (G367gat, keyinput26, G367gat_enc);
nand NAND2_96 (G368gat_enc, G43gat, G275gat);
xnor XNOR2_97 (G368gat, keyinput27, G368gat_enc);
nand NAND2_98 (G369gat_enc, G50gat, G275gat);
xor XOR2_99 (G369gat, keyinput28, G369gat_enc);
nand NAND2_100 (G370gat_enc, G57gat, G278gat);
xnor XNOR2_101 (G370gat, keyinput29, G370gat_enc);
nand NAND2_102 (G371gat_enc, G64gat, G278gat);
xor XOR2_103 (G371gat, keyinput30, G371gat_enc);
nand NAND2_104 (G372gat, G71gat, G281gat);
nand NAND2_105 (G373gat, G78gat, G281gat);
nand NAND2_106 (G374gat_enc, G85gat, G284gat);
xnor XNOR2_107 (G374gat, keyinput31, G374gat_enc);
nand NAND2_108 (G375gat, G92gat, G284gat);
nand NAND2_109 (G376gat, G99gat, G287gat);
nand NAND2_110 (G377gat, G106gat, G287gat);
nand NAND2_111 (G378gat, G113gat, G290gat);
nand NAND2_112 (G379gat, G120gat, G290gat);
nand NAND2_113 (G380gat, G127gat, G293gat);
nand NAND2_114 (G381gat, G134gat, G293gat);
nand NAND2_115 (G382gat, G141gat, G296gat);
nand NAND2_116 (G383gat, G148gat, G296gat);
nand NAND2_117 (G384gat, G155gat, G299gat);
nand NAND2_118 (G385gat, G162gat, G299gat);
nand NAND2_119 (G386gat, G169gat, G302gat);
nand NAND2_120 (G387gat, G176gat, G302gat);
nand NAND2_121 (G388gat, G183gat, G305gat);
nand NAND2_122 (G389gat, G190gat, G305gat);
nand NAND2_123 (G390gat, G197gat, G308gat);
nand NAND2_124 (G391gat, G204gat, G308gat);
nand NAND2_125 (G392gat, G211gat, G311gat);
nand NAND2_126 (G393gat, G218gat, G311gat);
nand NAND2_127 (G394gat, G1gat, G314gat);
nand NAND2_128 (G395gat, G29gat, G314gat);
nand NAND2_129 (G396gat, G57gat, G317gat);
nand NAND2_130 (G397gat, G85gat, G317gat);
nand NAND2_131 (G398gat, G8gat, G320gat);
nand NAND2_132 (G399gat, G36gat, G320gat);
nand NAND2_133 (G400gat, G64gat, G323gat);
nand NAND2_134 (G401gat, G92gat, G323gat);
nand NAND2_135 (G402gat, G15gat, G326gat);
nand NAND2_136 (G403gat, G43gat, G326gat);
nand NAND2_137 (G404gat, G71gat, G329gat);
nand NAND2_138 (G405gat, G99gat, G329gat);
nand NAND2_139 (G406gat, G22gat, G332gat);
nand NAND2_140 (G407gat, G50gat, G332gat);
nand NAND2_141 (G408gat, G78gat, G335gat);
nand NAND2_142 (G409gat, G106gat, G335gat);
nand NAND2_143 (G410gat, G113gat, G338gat);
nand NAND2_144 (G411gat, G141gat, G338gat);
nand NAND2_145 (G412gat, G169gat, G341gat);
nand NAND2_146 (G413gat, G197gat, G341gat);
nand NAND2_147 (G414gat, G120gat, G344gat);
nand NAND2_148 (G415gat, G148gat, G344gat);
nand NAND2_149 (G416gat, G176gat, G347gat);
nand NAND2_150 (G417gat, G204gat, G347gat);
nand NAND2_151 (G418gat, G127gat, G350gat);
nand NAND2_152 (G419gat, G155gat, G350gat);
nand NAND2_153 (G420gat, G183gat, G353gat);
nand NAND2_154 (G421gat, G211gat, G353gat);
nand NAND2_155 (G422gat, G134gat, G356gat);
nand NAND2_156 (G423gat, G162gat, G356gat);
nand NAND2_157 (G424gat, G190gat, G359gat);
nand NAND2_158 (G425gat, G218gat, G359gat);
nand NAND2_159 (G426gat, G362gat, G363gat);
nand NAND2_160 (G429gat, G364gat, G365gat);
nand NAND2_161 (G432gat, G366gat, G367gat);
nand NAND2_162 (G435gat, G368gat, G369gat);
nand NAND2_163 (G438gat, G370gat, G371gat);
nand NAND2_164 (G441gat, G372gat, G373gat);
nand NAND2_165 (G444gat, G374gat, G375gat);
nand NAND2_166 (G447gat, G376gat, G377gat);
nand NAND2_167 (G450gat, G378gat, G379gat);
nand NAND2_168 (G453gat, G380gat, G381gat);
nand NAND2_169 (G456gat, G382gat, G383gat);
nand NAND2_170 (G459gat, G384gat, G385gat);
nand NAND2_171 (G462gat, G386gat, G387gat);
nand NAND2_172 (G465gat, G388gat, G389gat);
nand NAND2_173 (G468gat, G390gat, G391gat);
nand NAND2_174 (G471gat, G392gat, G393gat);
nand NAND2_175 (G474gat, G394gat, G395gat);
nand NAND2_176 (G477gat, G396gat, G397gat);
nand NAND2_177 (G480gat, G398gat, G399gat);
nand NAND2_178 (G483gat, G400gat, G401gat);
nand NAND2_179 (G486gat, G402gat, G403gat);
nand NAND2_180 (G489gat, G404gat, G405gat);
nand NAND2_181 (G492gat, G406gat, G407gat);
nand NAND2_182 (G495gat, G408gat, G409gat);
nand NAND2_183 (G498gat, G410gat, G411gat);
nand NAND2_184 (G501gat, G412gat, G413gat);
nand NAND2_185 (G504gat, G414gat, G415gat);
nand NAND2_186 (G507gat, G416gat, G417gat);
nand NAND2_187 (G510gat, G418gat, G419gat);
nand NAND2_188 (G513gat, G420gat, G421gat);
nand NAND2_189 (G516gat, G422gat, G423gat);
nand NAND2_190 (G519gat, G424gat, G425gat);
nand NAND2_191 (G522gat, G426gat, G429gat);
nand NAND2_192 (G525gat, G432gat, G435gat);
nand NAND2_193 (G528gat, G438gat, G441gat);
nand NAND2_194 (G531gat, G444gat, G447gat);
nand NAND2_195 (G534gat, G450gat, G453gat);
nand NAND2_196 (G537gat, G456gat, G459gat);
nand NAND2_197 (G540gat, G462gat, G465gat);
nand NAND2_198 (G543gat, G468gat, G471gat);
nand NAND2_199 (G546gat, G474gat, G477gat);
nand NAND2_200 (G549gat, G480gat, G483gat);
nand NAND2_201 (G552gat, G486gat, G489gat);
nand NAND2_202 (G555gat, G492gat, G495gat);
nand NAND2_203 (G558gat, G498gat, G501gat);
nand NAND2_204 (G561gat, G504gat, G507gat);
nand NAND2_205 (G564gat, G510gat, G513gat);
nand NAND2_206 (G567gat, G516gat, G519gat);
nand NAND2_207 (G570gat, G426gat, G522gat);
nand NAND2_208 (G571gat, G429gat, G522gat);
nand NAND2_209 (G572gat, G432gat, G525gat);
nand NAND2_210 (G573gat, G435gat, G525gat);
nand NAND2_211 (G574gat, G438gat, G528gat);
nand NAND2_212 (G575gat, G441gat, G528gat);
nand NAND2_213 (G576gat, G444gat, G531gat);
nand NAND2_214 (G577gat, G447gat, G531gat);
nand NAND2_215 (G578gat, G450gat, G534gat);
nand NAND2_216 (G579gat, G453gat, G534gat);
nand NAND2_217 (G580gat, G456gat, G537gat);
nand NAND2_218 (G581gat, G459gat, G537gat);
nand NAND2_219 (G582gat, G462gat, G540gat);
nand NAND2_220 (G583gat, G465gat, G540gat);
nand NAND2_221 (G584gat, G468gat, G543gat);
nand NAND2_222 (G585gat, G471gat, G543gat);
nand NAND2_223 (G586gat, G474gat, G546gat);
nand NAND2_224 (G587gat, G477gat, G546gat);
nand NAND2_225 (G588gat, G480gat, G549gat);
nand NAND2_226 (G589gat, G483gat, G549gat);
nand NAND2_227 (G590gat, G486gat, G552gat);
nand NAND2_228 (G591gat, G489gat, G552gat);
nand NAND2_229 (G592gat, G492gat, G555gat);
nand NAND2_230 (G593gat, G495gat, G555gat);
nand NAND2_231 (G594gat, G498gat, G558gat);
nand NAND2_232 (G595gat, G501gat, G558gat);
nand NAND2_233 (G596gat, G504gat, G561gat);
nand NAND2_234 (G597gat, G507gat, G561gat);
nand NAND2_235 (G598gat, G510gat, G564gat);
nand NAND2_236 (G599gat, G513gat, G564gat);
nand NAND2_237 (G600gat, G516gat, G567gat);
nand NAND2_238 (G601gat, G519gat, G567gat);
nand NAND2_239 (G602gat, G570gat, G571gat);
nand NAND2_240 (G607gat, G572gat, G573gat);
nand NAND2_241 (G612gat, G574gat, G575gat);
nand NAND2_242 (G617gat, G576gat, G577gat);
nand NAND2_243 (G622gat, G578gat, G579gat);
nand NAND2_244 (G627gat, G580gat, G581gat);
nand NAND2_245 (G632gat, G582gat, G583gat);
nand NAND2_246 (G637gat, G584gat, G585gat);
nand NAND2_247 (G642gat, G586gat, G587gat);
nand NAND2_248 (G645gat, G588gat, G589gat);
nand NAND2_249 (G648gat, G590gat, G591gat);
nand NAND2_250 (G651gat, G592gat, G593gat);
nand NAND2_251 (G654gat, G594gat, G595gat);
nand NAND2_252 (G657gat, G596gat, G597gat);
nand NAND2_253 (G660gat, G598gat, G599gat);
nand NAND2_254 (G663gat, G600gat, G601gat);
nand NAND2_255 (G666gat, G602gat, G607gat);
nand NAND2_256 (G669gat, G612gat, G617gat);
nand NAND2_257 (G672gat, G602gat, G612gat);
nand NAND2_258 (G675gat, G607gat, G617gat);
nand NAND2_259 (G678gat, G622gat, G627gat);
nand NAND2_260 (G681gat, G632gat, G637gat);
nand NAND2_261 (G684gat, G622gat, G632gat);
nand NAND2_262 (G687gat, G627gat, G637gat);
nand NAND2_263 (G690gat, G602gat, G666gat);
nand NAND2_264 (G691gat, G607gat, G666gat);
nand NAND2_265 (G692gat, G612gat, G669gat);
nand NAND2_266 (G693gat, G617gat, G669gat);
nand NAND2_267 (G694gat, G602gat, G672gat);
nand NAND2_268 (G695gat, G612gat, G672gat);
nand NAND2_269 (G696gat, G607gat, G675gat);
nand NAND2_270 (G697gat, G617gat, G675gat);
nand NAND2_271 (G698gat, G622gat, G678gat);
nand NAND2_272 (G699gat, G627gat, G678gat);
nand NAND2_273 (G700gat, G632gat, G681gat);
nand NAND2_274 (G701gat, G637gat, G681gat);
nand NAND2_275 (G702gat, G622gat, G684gat);
nand NAND2_276 (G703gat, G632gat, G684gat);
nand NAND2_277 (G704gat, G627gat, G687gat);
nand NAND2_278 (G705gat, G637gat, G687gat);
nand NAND2_279 (G706gat, G690gat, G691gat);
nand NAND2_280 (G709gat, G692gat, G693gat);
nand NAND2_281 (G712gat, G694gat, G695gat);
nand NAND2_282 (G715gat, G696gat, G697gat);
nand NAND2_283 (G718gat, G698gat, G699gat);
nand NAND2_284 (G721gat, G700gat, G701gat);
nand NAND2_285 (G724gat, G702gat, G703gat);
nand NAND2_286 (G727gat, G704gat, G705gat);
nand NAND2_287 (G730gat, G242gat, G718gat);
nand NAND2_288 (G733gat, G245gat, G721gat);
nand NAND2_289 (G736gat, G248gat, G724gat);
nand NAND2_290 (G739gat, G251gat, G727gat);
nand NAND2_291 (G742gat, G254gat, G706gat);
nand NAND2_292 (G745gat, G257gat, G709gat);
nand NAND2_293 (G748gat, G260gat, G712gat);
nand NAND2_294 (G751gat, G263gat, G715gat);
nand NAND2_295 (G754gat, G242gat, G730gat);
nand NAND2_296 (G755gat, G718gat, G730gat);
nand NAND2_297 (G756gat, G245gat, G733gat);
nand NAND2_298 (G757gat, G721gat, G733gat);
nand NAND2_299 (G758gat, G248gat, G736gat);
nand NAND2_300 (G759gat, G724gat, G736gat);
nand NAND2_301 (G760gat, G251gat, G739gat);
nand NAND2_302 (G761gat, G727gat, G739gat);
nand NAND2_303 (G762gat, G254gat, G742gat);
nand NAND2_304 (G763gat, G706gat, G742gat);
nand NAND2_305 (G764gat, G257gat, G745gat);
nand NAND2_306 (G765gat, G709gat, G745gat);
nand NAND2_307 (G766gat, G260gat, G748gat);
nand NAND2_308 (G767gat, G712gat, G748gat);
nand NAND2_309 (G768gat, G263gat, G751gat);
nand NAND2_310 (G769gat, G715gat, G751gat);
nand NAND2_311 (G770gat, G754gat, G755gat);
nand NAND2_312 (G773gat, G756gat, G757gat);
nand NAND2_313 (G776gat, G758gat, G759gat);
nand NAND2_314 (G779gat, G760gat, G761gat);
nand NAND2_315 (G782gat, G762gat, G763gat);
nand NAND2_316 (G785gat, G764gat, G765gat);
nand NAND2_317 (G788gat, G766gat, G767gat);
nand NAND2_318 (G791gat, G768gat, G769gat);
nand NAND2_319 (G794gat, G642gat, G770gat);
nand NAND2_320 (G797gat, G645gat, G773gat);
nand NAND2_321 (G800gat, G648gat, G776gat);
nand NAND2_322 (G803gat, G651gat, G779gat);
nand NAND2_323 (G806gat, G654gat, G782gat);
nand NAND2_324 (G809gat, G657gat, G785gat);
nand NAND2_325 (G812gat, G660gat, G788gat);
nand NAND2_326 (G815gat, G663gat, G791gat);
nand NAND2_327 (G818gat, G642gat, G794gat);
nand NAND2_328 (G819gat, G770gat, G794gat);
nand NAND2_329 (G820gat, G645gat, G797gat);
nand NAND2_330 (G821gat, G773gat, G797gat);
nand NAND2_331 (G822gat, G648gat, G800gat);
nand NAND2_332 (G823gat, G776gat, G800gat);
nand NAND2_333 (G824gat, G651gat, G803gat);
nand NAND2_334 (G825gat, G779gat, G803gat);
nand NAND2_335 (G826gat, G654gat, G806gat);
nand NAND2_336 (G827gat, G782gat, G806gat);
nand NAND2_337 (G828gat, G657gat, G809gat);
nand NAND2_338 (G829gat, G785gat, G809gat);
nand NAND2_339 (G830gat, G660gat, G812gat);
nand NAND2_340 (G831gat, G788gat, G812gat);
nand NAND2_341 (G832gat, G663gat, G815gat);
nand NAND2_342 (G833gat, G791gat, G815gat);
nand NAND2_343 (G834gat, G818gat, G819gat);
nand NAND2_344 (G847gat, G820gat, G821gat);
nand NAND2_345 (G860gat, G822gat, G823gat);
nand NAND2_346 (G873gat, G824gat, G825gat);
nand NAND2_347 (G886gat, G828gat, G829gat);
nand NAND2_348 (G899gat, G832gat, G833gat);
nand NAND2_349 (G912gat, G830gat, G831gat);
nand NAND2_350 (G925gat, G826gat, G827gat);
not NOT1_351 (G938gat, G834gat);
not NOT1_352 (G939gat, G847gat);
not NOT1_353 (G940gat, G860gat);
not NOT1_354 (G941gat, G834gat);
not NOT1_355 (G942gat, G847gat);
not NOT1_356 (G943gat, G873gat);
not NOT1_357 (G944gat, G834gat);
not NOT1_358 (G945gat, G860gat);
not NOT1_359 (G946gat, G873gat);
not NOT1_360 (G947gat, G847gat);
not NOT1_361 (G948gat, G860gat);
not NOT1_362 (G949gat, G873gat);
not NOT1_363 (G950gat, G886gat);
not NOT1_364 (G951gat, G899gat);
not NOT1_365 (G952gat, G886gat);
not NOT1_366 (G953gat, G912gat);
not NOT1_367 (G954gat, G925gat);
not NOT1_368 (G955gat, G899gat);
not NOT1_369 (G956gat, G925gat);
not NOT1_370 (G957gat, G912gat);
not NOT1_371 (G958gat, G925gat);
not NOT1_372 (G959gat, G886gat);
not NOT1_373 (G960gat, G912gat);
not NOT1_374 (G961gat, G925gat);
not NOT1_375 (G962gat, G886gat);
not NOT1_376 (G963gat, G899gat);
not NOT1_377 (G964gat, G925gat);
not NOT1_378 (G965gat, G912gat);
not NOT1_379 (G966gat, G899gat);
not NOT1_380 (G967gat, G886gat);
not NOT1_381 (G968gat, G912gat);
not NOT1_382 (G969gat, G899gat);
not NOT1_383 (G970gat, G847gat);
not NOT1_384 (G971gat, G873gat);
not NOT1_385 (G972gat, G847gat);
not NOT1_386 (G973gat, G860gat);
not NOT1_387 (G974gat, G834gat);
not NOT1_388 (G975gat, G873gat);
not NOT1_389 (G976gat, G834gat);
not NOT1_390 (G977gat, G860gat);
and AND4_391 (G978gat, G938gat, G939gat, G940gat, G873gat);
and AND4_392 (G979gat, G941gat, G942gat, G860gat, G943gat);
and AND4_393 (G980gat, G944gat, G847gat, G945gat, G946gat);
and AND4_394 (G981gat, G834gat, G947gat, G948gat, G949gat);
and AND4_395 (G982gat, G958gat, G959gat, G960gat, G899gat);
and AND4_396 (G983gat, G961gat, G962gat, G912gat, G963gat);
and AND4_397 (G984gat, G964gat, G886gat, G965gat, G966gat);
and AND4_398 (G985gat, G925gat, G967gat, G968gat, G969gat);
or OR4_399 (G986gat, G978gat, G979gat, G980gat, G981gat);
or OR4_400 (G991gat, G982gat, G983gat, G984gat, G985gat);
and AND5_401 (G996gat, G925gat, G950gat, G912gat, G951gat, G986gat);
and AND5_402 (G1001gat, G925gat, G952gat, G953gat, G899gat, G986gat);
and AND5_403 (G1006gat, G954gat, G886gat, G912gat, G955gat, G986gat);
and AND5_404 (G1011gat, G956gat, G886gat, G957gat, G899gat, G986gat);
and AND5_405 (G1016gat, G834gat, G970gat, G860gat, G971gat, G991gat);
and AND5_406 (G1021gat, G834gat, G972gat, G973gat, G873gat, G991gat);
and AND5_407 (G1026gat, G974gat, G847gat, G860gat, G975gat, G991gat);
and AND5_408 (G1031gat, G976gat, G847gat, G977gat, G873gat, G991gat);
and AND2_409 (G1036gat, G834gat, G996gat);
and AND2_410 (G1039gat, G847gat, G996gat);
and AND2_411 (G1042gat, G860gat, G996gat);
and AND2_412 (G1045gat, G873gat, G996gat);
and AND2_413 (G1048gat, G834gat, G1001gat);
and AND2_414 (G1051gat, G847gat, G1001gat);
and AND2_415 (G1054gat, G860gat, G1001gat);
and AND2_416 (G1057gat, G873gat, G1001gat);
and AND2_417 (G1060gat, G834gat, G1006gat);
and AND2_418 (G1063gat, G847gat, G1006gat);
and AND2_419 (G1066gat, G860gat, G1006gat);
and AND2_420 (G1069gat, G873gat, G1006gat);
and AND2_421 (G1072gat, G834gat, G1011gat);
and AND2_422 (G1075gat, G847gat, G1011gat);
and AND2_423 (G1078gat, G860gat, G1011gat);
and AND2_424 (G1081gat, G873gat, G1011gat);
and AND2_425 (G1084gat, G925gat, G1016gat);
and AND2_426 (G1087gat, G886gat, G1016gat);
and AND2_427 (G1090gat, G912gat, G1016gat);
and AND2_428 (G1093gat, G899gat, G1016gat);
and AND2_429 (G1096gat, G925gat, G1021gat);
and AND2_430 (G1099gat, G886gat, G1021gat);
and AND2_431 (G1102gat, G912gat, G1021gat);
and AND2_432 (G1105gat, G899gat, G1021gat);
and AND2_433 (G1108gat, G925gat, G1026gat);
and AND2_434 (G1111gat, G886gat, G1026gat);
and AND2_435 (G1114gat, G912gat, G1026gat);
and AND2_436 (G1117gat, G899gat, G1026gat);
and AND2_437 (G1120gat, G925gat, G1031gat);
and AND2_438 (G1123gat, G886gat, G1031gat);
and AND2_439 (G1126gat, G912gat, G1031gat);
and AND2_440 (G1129gat, G899gat, G1031gat);
nand NAND2_441 (G1132gat, G1gat, G1036gat);
nand NAND2_442 (G1135gat, G8gat, G1039gat);
nand NAND2_443 (G1138gat, G15gat, G1042gat);
nand NAND2_444 (G1141gat, G22gat, G1045gat);
nand NAND2_445 (G1144gat, G29gat, G1048gat);
nand NAND2_446 (G1147gat, G36gat, G1051gat);
nand NAND2_447 (G1150gat, G43gat, G1054gat);
nand NAND2_448 (G1153gat, G50gat, G1057gat);
nand NAND2_449 (G1156gat, G57gat, G1060gat);
nand NAND2_450 (G1159gat, G64gat, G1063gat);
nand NAND2_451 (G1162gat, G71gat, G1066gat);
nand NAND2_452 (G1165gat, G78gat, G1069gat);
nand NAND2_453 (G1168gat, G85gat, G1072gat);
nand NAND2_454 (G1171gat, G92gat, G1075gat);
nand NAND2_455 (G1174gat, G99gat, G1078gat);
nand NAND2_456 (G1177gat, G106gat, G1081gat);
nand NAND2_457 (G1180gat, G113gat, G1084gat);
nand NAND2_458 (G1183gat, G120gat, G1087gat);
nand NAND2_459 (G1186gat, G127gat, G1090gat);
nand NAND2_460 (G1189gat, G134gat, G1093gat);
nand NAND2_461 (G1192gat, G141gat, G1096gat);
nand NAND2_462 (G1195gat, G148gat, G1099gat);
nand NAND2_463 (G1198gat, G155gat, G1102gat);
nand NAND2_464 (G1201gat, G162gat, G1105gat);
nand NAND2_465 (G1204gat, G169gat, G1108gat);
nand NAND2_466 (G1207gat, G176gat, G1111gat);
nand NAND2_467 (G1210gat, G183gat, G1114gat);
nand NAND2_468 (G1213gat, G190gat, G1117gat);
nand NAND2_469 (G1216gat, G197gat, G1120gat);
nand NAND2_470 (G1219gat, G204gat, G1123gat);
nand NAND2_471 (G1222gat, G211gat, G1126gat);
nand NAND2_472 (G1225gat, G218gat, G1129gat);
nand NAND2_473 (G1228gat, G1gat, G1132gat);
nand NAND2_474 (G1229gat, G1036gat, G1132gat);
nand NAND2_475 (G1230gat, G8gat, G1135gat);
nand NAND2_476 (G1231gat, G1039gat, G1135gat);
nand NAND2_477 (G1232gat, G15gat, G1138gat);
nand NAND2_478 (G1233gat, G1042gat, G1138gat);
nand NAND2_479 (G1234gat, G22gat, G1141gat);
nand NAND2_480 (G1235gat, G1045gat, G1141gat);
nand NAND2_481 (G1236gat, G29gat, G1144gat);
nand NAND2_482 (G1237gat, G1048gat, G1144gat);
nand NAND2_483 (G1238gat, G36gat, G1147gat);
nand NAND2_484 (G1239gat, G1051gat, G1147gat);
nand NAND2_485 (G1240gat, G43gat, G1150gat);
nand NAND2_486 (G1241gat, G1054gat, G1150gat);
nand NAND2_487 (G1242gat, G50gat, G1153gat);
nand NAND2_488 (G1243gat, G1057gat, G1153gat);
nand NAND2_489 (G1244gat, G57gat, G1156gat);
nand NAND2_490 (G1245gat, G1060gat, G1156gat);
nand NAND2_491 (G1246gat, G64gat, G1159gat);
nand NAND2_492 (G1247gat, G1063gat, G1159gat);
nand NAND2_493 (G1248gat, G71gat, G1162gat);
nand NAND2_494 (G1249gat, G1066gat, G1162gat);
nand NAND2_495 (G1250gat, G78gat, G1165gat);
nand NAND2_496 (G1251gat, G1069gat, G1165gat);
nand NAND2_497 (G1252gat, G85gat, G1168gat);
nand NAND2_498 (G1253gat, G1072gat, G1168gat);
nand NAND2_499 (G1254gat, G92gat, G1171gat);
nand NAND2_500 (G1255gat, G1075gat, G1171gat);
nand NAND2_501 (G1256gat, G99gat, G1174gat);
nand NAND2_502 (G1257gat, G1078gat, G1174gat);
nand NAND2_503 (G1258gat, G106gat, G1177gat);
nand NAND2_504 (G1259gat, G1081gat, G1177gat);
nand NAND2_505 (G1260gat, G113gat, G1180gat);
nand NAND2_506 (G1261gat, G1084gat, G1180gat);
nand NAND2_507 (G1262gat, G120gat, G1183gat);
nand NAND2_508 (G1263gat, G1087gat, G1183gat);
nand NAND2_509 (G1264gat, G127gat, G1186gat);
nand NAND2_510 (G1265gat, G1090gat, G1186gat);
nand NAND2_511 (G1266gat, G134gat, G1189gat);
nand NAND2_512 (G1267gat, G1093gat, G1189gat);
nand NAND2_513 (G1268gat, G141gat, G1192gat);
nand NAND2_514 (G1269gat, G1096gat, G1192gat);
nand NAND2_515 (G1270gat, G148gat, G1195gat);
nand NAND2_516 (G1271gat, G1099gat, G1195gat);
nand NAND2_517 (G1272gat, G155gat, G1198gat);
nand NAND2_518 (G1273gat, G1102gat, G1198gat);
nand NAND2_519 (G1274gat, G162gat, G1201gat);
nand NAND2_520 (G1275gat, G1105gat, G1201gat);
nand NAND2_521 (G1276gat, G169gat, G1204gat);
nand NAND2_522 (G1277gat, G1108gat, G1204gat);
nand NAND2_523 (G1278gat, G176gat, G1207gat);
nand NAND2_524 (G1279gat, G1111gat, G1207gat);
nand NAND2_525 (G1280gat, G183gat, G1210gat);
nand NAND2_526 (G1281gat, G1114gat, G1210gat);
nand NAND2_527 (G1282gat, G190gat, G1213gat);
nand NAND2_528 (G1283gat, G1117gat, G1213gat);
nand NAND2_529 (G1284gat, G197gat, G1216gat);
nand NAND2_530 (G1285gat, G1120gat, G1216gat);
nand NAND2_531 (G1286gat, G204gat, G1219gat);
nand NAND2_532 (G1287gat, G1123gat, G1219gat);
nand NAND2_533 (G1288gat, G211gat, G1222gat);
nand NAND2_534 (G1289gat, G1126gat, G1222gat);
nand NAND2_535 (G1290gat, G218gat, G1225gat);
nand NAND2_536 (G1291gat, G1129gat, G1225gat);
nand NAND2_537 (G1292gat, G1228gat, G1229gat);
nand NAND2_538 (G1293gat, G1230gat, G1231gat);
nand NAND2_539 (G1294gat, G1232gat, G1233gat);
nand NAND2_540 (G1295gat, G1234gat, G1235gat);
nand NAND2_541 (G1296gat, G1236gat, G1237gat);
nand NAND2_542 (G1297gat, G1238gat, G1239gat);
nand NAND2_543 (G1298gat, G1240gat, G1241gat);
nand NAND2_544 (G1299gat, G1242gat, G1243gat);
nand NAND2_545 (G1300gat, G1244gat, G1245gat);
nand NAND2_546 (G1301gat, G1246gat, G1247gat);
nand NAND2_547 (G1302gat, G1248gat, G1249gat);
nand NAND2_548 (G1303gat, G1250gat, G1251gat);
nand NAND2_549 (G1304gat, G1252gat, G1253gat);
nand NAND2_550 (G1305gat, G1254gat, G1255gat);
nand NAND2_551 (G1306gat, G1256gat, G1257gat);
nand NAND2_552 (G1307gat, G1258gat, G1259gat);
nand NAND2_553 (G1308gat, G1260gat, G1261gat);
nand NAND2_554 (G1309gat, G1262gat, G1263gat);
nand NAND2_555 (G1310gat, G1264gat, G1265gat);
nand NAND2_556 (G1311gat, G1266gat, G1267gat);
nand NAND2_557 (G1312gat, G1268gat, G1269gat);
nand NAND2_558 (G1313gat, G1270gat, G1271gat);
nand NAND2_559 (G1314gat, G1272gat, G1273gat);
nand NAND2_560 (G1315gat, G1274gat, G1275gat);
nand NAND2_561 (G1316gat, G1276gat, G1277gat);
nand NAND2_562 (G1317gat, G1278gat, G1279gat);
nand NAND2_563 (G1318gat, G1280gat, G1281gat);
nand NAND2_564 (G1319gat, G1282gat, G1283gat);
nand NAND2_565 (G1320gat, G1284gat, G1285gat);
nand NAND2_566 (G1321gat, G1286gat, G1287gat);
nand NAND2_567 (G1322gat, G1288gat, G1289gat);
nand NAND2_568 (G1323gat, G1290gat, G1291gat);

endmodule