module DFF(Q, clk, D);
input D;
input clk;
output Q;
always @(clk)
begin
  Q <= D;
end
endmodule


module c432_libar_16k(G1gat,G4gat,G8gat,G11gat,G14gat,G17gat,G21gat,G24gat,G27gat,G30gat,G34gat,G37gat,G40gat,G43gat,G47gat,G50gat,G53gat,G56gat,G60gat,G63gat,G66gat,G69gat,G73gat,G76gat,G79gat,G82gat,G86gat,G89gat,G92gat,G95gat,G99gat,G102gat,G105gat,G108gat,G112gat,G115gat,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15,G223gat,G329gat,G370gat,G421gat,G430gat,G431gat,G432gat);

input G1gat,G4gat,G8gat,G11gat,G14gat,G17gat,G21gat,G24gat,G27gat,G30gat,G34gat,G37gat,G40gat,G43gat,G47gat,G50gat,G53gat,G56gat,G60gat,G63gat,G66gat,G69gat,G73gat,G76gat,G79gat,G82gat,G86gat,G89gat,G92gat,G95gat,G99gat,G102gat,G105gat,G108gat,G112gat,G115gat,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15;
output G223gat,G329gat,G370gat,G421gat,G430gat,G431gat,G432gat;
wire G118gat,G119gat,G122gat_enc,G122gat,G123gat,G126gat,G127gat_enc,G127gat,G130gat_enc,G130gat,G131gat_enc,CLK8,LIBAR8,G131gat,G134gat_enc,G134gat,G135gat,G138gat,G139gat_enc,G139gat,G142gat_enc,G142gat,G143gat_enc,G143gat,G146gat,G147gat_enc,G147gat,G150gat_enc,CLK7,LIBAR7,G150gat,G151gat_enc,CLK6,LIBAR6,G151gat,G154gat_enc,CLK5,LIBAR5,G154gat,G157gat_enc,CLK4,LIBAR4,G157gat,G158gat_enc,CLK3,LIBAR3,G158gat,G159gat_enc,CLK2,LIBAR2,G159gat,G162gat_enc,CLK1,LIBAR1,G162gat,G165gat,G168gat,G171gat,G174gat,G177gat,G180gat,G183gat,G184gat,G185gat,G186gat,G187gat,G188gat,G189gat,G190gat,G191gat,G192gat,G193gat,G194gat,G195gat,G196gat,G197gat,G198gat,G1980gat,G1981gat,G199gat,G203gat,G213gat,G224gat,G227gat,G230gat,G233gat,G236gat,G239gat,G242gat,G243gat,G246gat,G247gat,G250gat,G251gat,G254gat,G255gat,G256gat,G257gat,G258gat,G259gat,G260gat,G263gat,G264gat,G267gat,G270gat,G273gat,G276gat,G279gat,G282gat,G285gat,G288gat,G289gat,G290gat,G291gat,G292gat,G293gat,G294gat,G295gat,G2950gat,G2951gat,G296gat,G300gat,G301gat,G302gat,G303gat,G304gat,G305gat,G306gat,G307gat,G308gat,G309gat,G319gat,G330gat,G331gat,G332gat,G333gat,G334gat,G335gat,G336gat,G337gat,G338gat,G339gat,G340gat,G341gat,G342gat,G343gat,G344gat,G345gat,G346gat,G347gat,G348gat,G349gat,G350gat,G351gat,G352gat,G353gat,G354gat,G355gat,G356gat,G3560gat,G3561gat,G357gat,G360gat,G371gat,G372gat,G373gat,G374gat,G375gat,G376gat,G377gat,G378gat,G379gat,G380gat,G381gat,G386gat,G393gat,G399gat,G404gat,G407gat,G411gat,G414gat,G415gat,G4150gat,G4151gat,G416gat,G417gat,G418gat,G419gat,G420gat,G422gat,G425gat,G428gat,G429gat;

not NOT1_1 (G118gat, G1gat);
not NOT1_2 (G119gat, G4gat);
not NOT1_3 (G122gat_enc, G11gat);
xnor XNOR2_4 (G122gat, keyinput0, G122gat_enc);
not NOT1_5 (G123gat, G17gat);
not NOT1_6 (G126gat, G24gat);
not NOT1_7 (G127gat_enc, G30gat);
xnor XNOR2_8 (G127gat, keyinput1, G127gat_enc);
not NOT1_9 (G130gat_enc, G37gat);
xor XOR2_10 (G130gat, keyinput2, G130gat_enc);
not NOT1_11 (G131gat_enc, G43gat);
nor NOR2_12 (CLK8, G131gat_enc, G130gat);
dff DFF2_13 (LIBAR8, CLK8, keyinput3);
xor XOR2_14 (G131gat, LIBAR8, G131gat_enc);
not NOT1_15 (G134gat_enc, G50gat);
xor XOR2_16 (G134gat, keyinput4, G134gat_enc);
not NOT1_17 (G135gat, G56gat);
not NOT1_18 (G138gat, G63gat);
not NOT1_19 (G139gat_enc, G69gat);
xnor XNOR2_20 (G139gat, keyinput5, G139gat_enc);
not NOT1_21 (G142gat_enc, G76gat);
xnor XNOR2_22 (G142gat, keyinput6, G142gat_enc);
not NOT1_23 (G143gat_enc, G82gat);
xor XOR2_24 (G143gat, keyinput7, G143gat_enc);
not NOT1_25 (G146gat, G89gat);
not NOT1_26 (G147gat_enc, G95gat);
xnor XNOR2_27 (G147gat, keyinput8, G147gat_enc);
not NOT1_28 (G150gat_enc, G102gat);
nor NOR2_29 (CLK7, G150gat_enc, G147gat);
dff DFF2_30 (LIBAR7, CLK7, keyinput9);
xor XOR2_31 (G150gat, LIBAR7, G150gat_enc);
not NOT1_32 (G151gat_enc, G108gat);
nor NOR2_33 (CLK6, G151gat_enc, G150gat);
dff DFF2_34 (LIBAR6, CLK6, keyinput10);
xnor XNOR2_35 (G151gat, LIBAR6, G151gat_enc);
nand NAND2_36 (G154gat_enc, G118gat, G4gat);
nor NOR2_37 (CLK5, G154gat_enc, G151gat);
dff DFF2_38 (LIBAR5, CLK5, keyinput11);
xor XOR2_39 (G154gat, LIBAR5, G154gat_enc);
nor NOR2_40 (G157gat_enc, G8gat, G119gat);
nor NOR2_41 (CLK4, G157gat_enc, G154gat);
dff DFF2_42 (LIBAR4, CLK4, keyinput12);
xnor XNOR2_43 (G157gat, LIBAR4, G157gat_enc);
nor NOR2_44 (G158gat_enc, G14gat, G119gat);
nor NOR2_45 (CLK3, G158gat_enc, G157gat);
dff DFF2_46 (LIBAR3, CLK3, keyinput13);
xnor XNOR2_47 (G158gat, LIBAR3, G158gat_enc);
nand NAND2_48 (G159gat_enc, G122gat, G17gat);
nor NOR2_49 (CLK2, G159gat_enc, G158gat);
dff DFF2_50 (LIBAR2, CLK2, keyinput14);
xor XOR2_51 (G159gat, LIBAR2, G159gat_enc);
nand NAND2_52 (G162gat_enc, G126gat, G30gat);
nor NOR2_53 (CLK1, G162gat_enc, G159gat);
dff DFF2_54 (LIBAR1, CLK1, keyinput15);
xor XOR2_55 (G162gat, LIBAR1, G162gat_enc);
nand NAND2_56 (G165gat, G130gat, G43gat);
nand NAND2_57 (G168gat, G134gat, G56gat);
nand NAND2_58 (G171gat, G138gat, G69gat);
nand NAND2_59 (G174gat, G142gat, G82gat);
nand NAND2_60 (G177gat, G146gat, G95gat);
nand NAND2_61 (G180gat, G150gat, G108gat);
nor NOR2_62 (G183gat, G21gat, G123gat);
nor NOR2_63 (G184gat, G27gat, G123gat);
nor NOR2_64 (G185gat, G34gat, G127gat);
nor NOR2_65 (G186gat, G40gat, G127gat);
nor NOR2_66 (G187gat, G47gat, G131gat);
nor NOR2_67 (G188gat, G53gat, G131gat);
nor NOR2_68 (G189gat, G60gat, G135gat);
nor NOR2_69 (G190gat, G66gat, G135gat);
nor NOR2_70 (G191gat, G73gat, G139gat);
nor NOR2_71 (G192gat, G79gat, G139gat);
nor NOR2_72 (G193gat, G86gat, G143gat);
nor NOR2_73 (G194gat, G92gat, G143gat);
nor NOR2_74 (G195gat, G99gat, G147gat);
nor NOR2_75 (G196gat, G105gat, G147gat);
nor NOR2_76 (G197gat, G112gat, G151gat);
nor NOR2_77 (G198gat, G115gat, G151gat);
and AND4_78 (G1980gat, G154gat, G159gat, G162gat, G165gat);
and AND5_79 (G1981gat, G168gat, G171gat, G174gat, G177gat, G180gat);
and AND2_80 (G199gat, G1980gat, G1981gat);
not NOT1_81 (G203gat, G199gat);
not NOT1_82 (G213gat, G199gat);
not NOT1_83 (G223gat, G199gat);
xor XOR2_84 (G224gat, G203gat, G154gat);
xor XOR2_85 (G227gat, G203gat, G159gat);
xor XOR2_86 (G230gat, G203gat, G162gat);
xor XOR2_87 (G233gat, G203gat, G165gat);
xor XOR2_88 (G236gat, G203gat, G168gat);
xor XOR2_89 (G239gat, G203gat, G171gat);
nand NAND2_90 (G242gat, G1gat, G213gat);
xor XOR2_91 (G243gat, G203gat, G174gat);
nand NAND2_92 (G246gat, G213gat, G11gat);
xor XOR2_93 (G247gat, G203gat, G177gat);
nand NAND2_94 (G250gat, G213gat, G24gat);
xor XOR2_95 (G251gat, G203gat, G180gat);
nand NAND2_96 (G254gat, G213gat, G37gat);
nand NAND2_97 (G255gat, G213gat, G50gat);
nand NAND2_98 (G256gat, G213gat, G63gat);
nand NAND2_99 (G257gat, G213gat, G76gat);
nand NAND2_100 (G258gat, G213gat, G89gat);
nand NAND2_101 (G259gat, G213gat, G102gat);
nand NAND2_102 (G260gat, G224gat, G157gat);
nand NAND2_103 (G263gat, G224gat, G158gat);
nand NAND2_104 (G264gat, G227gat, G183gat);
nand NAND2_105 (G267gat, G230gat, G185gat);
nand NAND2_106 (G270gat, G233gat, G187gat);
nand NAND2_107 (G273gat, G236gat, G189gat);
nand NAND2_108 (G276gat, G239gat, G191gat);
nand NAND2_109 (G279gat, G243gat, G193gat);
nand NAND2_110 (G282gat, G247gat, G195gat);
nand NAND2_111 (G285gat, G251gat, G197gat);
nand NAND2_112 (G288gat, G227gat, G184gat);
nand NAND2_113 (G289gat, G230gat, G186gat);
nand NAND2_114 (G290gat, G233gat, G188gat);
nand NAND2_115 (G291gat, G236gat, G190gat);
nand NAND2_116 (G292gat, G239gat, G192gat);
nand NAND2_117 (G293gat, G243gat, G194gat);
nand NAND2_118 (G294gat, G247gat, G196gat);
nand NAND2_119 (G295gat, G251gat, G198gat);
and AND4_120 (G2950gat, G260gat, G264gat, G267gat, G270gat);
and AND5_121 (G2951gat, G273gat, G276gat, G279gat, G282gat, G285gat);
and AND2_122 (G296gat, G2950gat, G2951gat);
not NOT1_123 (G300gat, G263gat);
not NOT1_124 (G301gat, G288gat);
not NOT1_125 (G302gat, G289gat);
not NOT1_126 (G303gat, G290gat);
not NOT1_127 (G304gat, G291gat);
not NOT1_128 (G305gat, G292gat);
not NOT1_129 (G306gat, G293gat);
not NOT1_130 (G307gat, G294gat);
not NOT1_131 (G308gat, G295gat);
not NOT1_132 (G309gat, G296gat);
not NOT1_133 (G319gat, G296gat);
not NOT1_134 (G329gat, G296gat);
xor XOR2_135 (G330gat, G309gat, G260gat);
xor XOR2_136 (G331gat, G309gat, G264gat);
xor XOR2_137 (G332gat, G309gat, G267gat);
xor XOR2_138 (G333gat, G309gat, G270gat);
nand NAND2_139 (G334gat, G8gat, G319gat);
xor XOR2_140 (G335gat, G309gat, G273gat);
nand NAND2_141 (G336gat, G319gat, G21gat);
xor XOR2_142 (G337gat, G309gat, G276gat);
nand NAND2_143 (G338gat, G319gat, G34gat);
xor XOR2_144 (G339gat, G309gat, G279gat);
nand NAND2_145 (G340gat, G319gat, G47gat);
xor XOR2_146 (G341gat, G309gat, G282gat);
nand NAND2_147 (G342gat, G319gat, G60gat);
xor XOR2_148 (G343gat, G309gat, G285gat);
nand NAND2_149 (G344gat, G319gat, G73gat);
nand NAND2_150 (G345gat, G319gat, G86gat);
nand NAND2_151 (G346gat, G319gat, G99gat);
nand NAND2_152 (G347gat, G319gat, G112gat);
nand NAND2_153 (G348gat, G330gat, G300gat);
nand NAND2_154 (G349gat, G331gat, G301gat);
nand NAND2_155 (G350gat, G332gat, G302gat);
nand NAND2_156 (G351gat, G333gat, G303gat);
nand NAND2_157 (G352gat, G335gat, G304gat);
nand NAND2_158 (G353gat, G337gat, G305gat);
nand NAND2_159 (G354gat, G339gat, G306gat);
nand NAND2_160 (G355gat, G341gat, G307gat);
nand NAND2_161 (G356gat, G343gat, G308gat);
and AND4_162 (G3560gat, G348gat, G349gat, G350gat, G351gat);
and AND5_163 (G3561gat, G352gat, G353gat, G354gat, G355gat, G356gat);
and AND2_164 (G357gat, G3560gat, G3561gat);
not NOT1_165 (G360gat, G357gat);
not NOT1_166 (G370gat, G357gat);
nand NAND2_167 (G371gat, G14gat, G360gat);
nand NAND2_168 (G372gat, G360gat, G27gat);
nand NAND2_169 (G373gat, G360gat, G40gat);
nand NAND2_170 (G374gat, G360gat, G53gat);
nand NAND2_171 (G375gat, G360gat, G66gat);
nand NAND2_172 (G376gat, G360gat, G79gat);
nand NAND2_173 (G377gat, G360gat, G92gat);
nand NAND2_174 (G378gat, G360gat, G105gat);
nand NAND2_175 (G379gat, G360gat, G115gat);
nand NAND4_176 (G380gat, G4gat, G242gat, G334gat, G371gat);
nand NAND4_177 (G381gat, G246gat, G336gat, G372gat, G17gat);
nand NAND4_178 (G386gat, G250gat, G338gat, G373gat, G30gat);
nand NAND4_179 (G393gat, G254gat, G340gat, G374gat, G43gat);
nand NAND4_180 (G399gat, G255gat, G342gat, G375gat, G56gat);
nand NAND4_181 (G404gat, G256gat, G344gat, G376gat, G69gat);
nand NAND4_182 (G407gat, G257gat, G345gat, G377gat, G82gat);
nand NAND4_183 (G411gat, G258gat, G346gat, G378gat, G95gat);
nand NAND4_184 (G414gat, G259gat, G347gat, G379gat, G108gat);
not NOT1_185 (G415gat, G380gat);
and AND4_186 (G4150gat, G381gat, G386gat, G393gat, G399gat);
and AND4_187 (G4151gat, G404gat, G407gat, G411gat, G414gat);
and AND2_188 (G416gat, G4150gat, G4151gat);
not NOT1_189 (G417gat, G393gat);
not NOT1_190 (G418gat, G404gat);
not NOT1_191 (G419gat, G407gat);
not NOT1_192 (G420gat, G411gat);
nor NOR2_193 (G421gat, G415gat, G416gat);
nand NAND2_194 (G422gat, G386gat, G417gat);
nand NAND4_195 (G425gat, G386gat, G393gat, G418gat, G399gat);
nand NAND3_196 (G428gat, G399gat, G393gat, G419gat);
nand NAND4_197 (G429gat, G386gat, G393gat, G407gat, G420gat);
nand NAND4_198 (G430gat, G381gat, G386gat, G422gat, G399gat);
nand NAND4_199 (G431gat, G381gat, G386gat, G425gat, G428gat);
nand NAND4_200 (G432gat, G381gat, G422gat, G425gat, G429gat);

endmodule