module DFF(Q, clk, D);
input D;
input clk;
output Q;
always @(clk)
begin
  Q <= D;
end
endmodule


module c6288_libar_16k(G1gat,G18gat,G35gat,G52gat,G69gat,G86gat,G103gat,G120gat,G137gat,G154gat,G171gat,G188gat,G205gat,G222gat,G239gat,G256gat,G273gat,G290gat,G307gat,G324gat,G341gat,G358gat,G375gat,G392gat,G409gat,G426gat,G443gat,G460gat,G477gat,G494gat,G511gat,G528gat,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15,G545gat,G1581gat,G1901gat,G2223gat,G2548gat,G2877gat,G3211gat,G3552gat,G3895gat,G4241gat,G4591gat,G4946gat,G5308gat,G5672gat,G5971gat,G6123gat,G6150gat,G6160gat,G6170gat,G6180gat,G6190gat,G6200gat,G6210gat,G6220gat,G6230gat,G6240gat,G6250gat,G6260gat,G6270gat,G6280gat,G6287gat,G6288gat);

input G1gat,G18gat,G35gat,G52gat,G69gat,G86gat,G103gat,G120gat,G137gat,G154gat,G171gat,G188gat,G205gat,G222gat,G239gat,G256gat,G273gat,G290gat,G307gat,G324gat,G341gat,G358gat,G375gat,G392gat,G409gat,G426gat,G443gat,G460gat,G477gat,G494gat,G511gat,G528gat,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15;
output G545gat,G1581gat,G1901gat,G2223gat,G2548gat,G2877gat,G3211gat,G3552gat,G3895gat,G4241gat,G4591gat,G4946gat,G5308gat,G5672gat,G5971gat,G6123gat,G6150gat,G6160gat,G6170gat,G6180gat,G6190gat,G6200gat,G6210gat,G6220gat,G6230gat,G6240gat,G6250gat,G6260gat,G6270gat,G6280gat,G6287gat,G6288gat;
wire G546gat,G549gat_enc,G549gat,G552gat,G555gat_enc,G555gat,G558gat_enc,CLK8,LIBAR8,G558gat,G561gat_enc,G561gat,G564gat_enc,G564gat,G567gat,G570gat_enc,G570gat,G573gat_enc,G573gat,G576gat_enc,G576gat,G579gat_enc,CLK7,LIBAR7,G579gat,G582gat_enc,G582gat,G585gat,G588gat,G591gat_enc,CLK6,LIBAR6,G591gat,G594gat_enc,CLK5,LIBAR5,G594gat,G597gat_enc,CLK4,LIBAR4,G597gat,G600gat,G603gat,G606gat_enc,CLK3,LIBAR3,G606gat,G609gat_enc,CLK2,LIBAR2,G609gat,G612gat_enc,CLK1,LIBAR1,G612gat,G615gat,G618gat,G621gat,G624gat,G627gat,G630gat,G633gat,G636gat,G639gat,G642gat,G645gat,G648gat,G651gat,G654gat,G657gat,G660gat,G663gat,G666gat,G669gat,G672gat,G675gat,G678gat,G681gat,G684gat,G687gat,G690gat,G693gat,G696gat,G699gat,G702gat,G705gat,G708gat,G711gat,G714gat,G717gat,G720gat,G723gat,G726gat,G729gat,G732gat,G735gat,G738gat,G741gat,G744gat,G747gat,G750gat,G753gat,G756gat,G759gat,G762gat,G765gat,G768gat,G771gat,G774gat,G777gat,G780gat,G783gat,G786gat,G789gat,G792gat,G795gat,G798gat,G801gat,G804gat,G807gat,G810gat,G813gat,G816gat,G819gat,G822gat,G825gat,G828gat,G831gat,G834gat,G837gat,G840gat,G843gat,G846gat,G849gat,G852gat,G855gat,G858gat,G861gat,G864gat,G867gat,G870gat,G873gat,G876gat,G879gat,G882gat,G885gat,G888gat,G891gat,G894gat,G897gat,G900gat,G903gat,G906gat,G909gat,G912gat,G915gat,G918gat,G921gat,G924gat,G927gat,G930gat,G933gat,G936gat,G939gat,G942gat,G945gat,G948gat,G951gat,G954gat,G957gat,G960gat,G963gat,G966gat,G969gat,G972gat,G975gat,G978gat,G981gat,G984gat,G987gat,G990gat,G993gat,G996gat,G999gat,G1002gat,G1005gat,G1008gat,G1011gat,G1014gat,G1017gat,G1020gat,G1023gat,G1026gat,G1029gat,G1032gat,G1035gat,G1038gat,G1041gat,G1044gat,G1047gat,G1050gat,G1053gat,G1056gat,G1059gat,G1062gat,G1065gat,G1068gat,G1071gat,G1074gat,G1077gat,G1080gat,G1083gat,G1086gat,G1089gat,G1092gat,G1095gat,G1098gat,G1101gat,G1104gat,G1107gat,G1110gat,G1113gat,G1116gat,G1119gat,G1122gat,G1125gat,G1128gat,G1131gat,G1134gat,G1137gat,G1140gat,G1143gat,G1146gat,G1149gat,G1152gat,G1155gat,G1158gat,G1161gat,G1164gat,G1167gat,G1170gat,G1173gat,G1176gat,G1179gat,G1182gat,G1185gat,G1188gat,G1191gat,G1194gat,G1197gat,G1200gat,G1203gat,G1206gat,G1209gat,G1212gat,G1215gat,G1218gat,G1221gat,G1224gat,G1227gat,G1230gat,G1233gat,G1236gat,G1239gat,G1242gat,G1245gat,G1248gat,G1251gat,G1254gat,G1257gat,G1260gat,G1263gat,G1266gat,G1269gat,G1272gat,G1275gat,G1278gat,G1281gat,G1284gat,G1287gat,G1290gat,G1293gat,G1296gat,G1299gat,G1302gat,G1305gat,G1308gat,G1311gat,G1315gat,G1319gat,G1323gat,G1327gat,G1331gat,G1335gat,G1339gat,G1343gat,G1347gat,G1351gat,G1355gat,G1359gat,G1363gat,G1367gat,G1371gat,G1372gat,G1373gat,G1374gat,G1375gat,G1376gat,G1377gat,G1378gat,G1379gat,G1380gat,G1381gat,G1382gat,G1383gat,G1384gat,G1385gat,G1386gat,G1387gat,G1388gat,G1389gat,G1390gat,G1391gat,G1392gat,G1393gat,G1394gat,G1395gat,G1396gat,G1397gat,G1398gat,G1399gat,G1400gat,G1401gat,G1404gat,G1407gat,G1410gat,G1413gat,G1416gat,G1419gat,G1422gat,G1425gat,G1428gat,G1431gat,G1434gat,G1437gat,G1440gat,G1443gat,G1446gat,G1450gat,G1454gat,G1458gat,G1462gat,G1466gat,G1470gat,G1474gat,G1478gat,G1482gat,G1486gat,G1490gat,G1494gat,G1498gat,G1502gat,G1506gat,G1507gat,G1508gat,G1511gat,G1512gat,G1513gat,G1516gat,G1517gat,G1518gat,G1521gat,G1522gat,G1523gat,G1526gat,G1527gat,G1528gat,G1531gat,G1532gat,G1533gat,G1536gat,G1537gat,G1538gat,G1541gat,G1542gat,G1543gat,G1546gat,G1547gat,G1548gat,G1551gat,G1552gat,G1553gat,G1556gat,G1557gat,G1558gat,G1561gat,G1562gat,G1563gat,G1566gat,G1567gat,G1568gat,G1571gat,G1572gat,G1573gat,G1576gat,G1577gat,G1578gat,G1582gat,G1585gat,G1588gat,G1591gat,G1594gat,G1597gat,G1600gat,G1603gat,G1606gat,G1609gat,G1612gat,G1615gat,G1618gat,G1621gat,G1624gat,G1628gat,G1632gat,G1636gat,G1640gat,G1644gat,G1648gat,G1652gat,G1656gat,G1660gat,G1664gat,G1668gat,G1672gat,G1676gat,G1680gat,G1684gat,G1685gat,G1686gat,G1687gat,G1688gat,G1689gat,G1690gat,G1691gat,G1692gat,G1693gat,G1694gat,G1695gat,G1696gat,G1697gat,G1698gat,G1699gat,G1700gat,G1701gat,G1702gat,G1703gat,G1704gat,G1705gat,G1706gat,G1707gat,G1708gat,G1709gat,G1710gat,G1711gat,G1712gat,G1713gat,G1714gat,G1717gat,G1720gat,G1723gat,G1726gat,G1729gat,G1732gat,G1735gat,G1738gat,G1741gat,G1744gat,G1747gat,G1750gat,G1753gat,G1756gat,G1759gat,G1763gat,G1767gat,G1771gat,G1775gat,G1779gat,G1783gat,G1787gat,G1791gat,G1795gat,G1799gat,G1803gat,G1807gat,G1811gat,G1815gat,G1819gat,G1820gat,G1821gat,G1824gat,G1825gat,G1826gat,G1829gat,G1830gat,G1831gat,G1834gat,G1835gat,G1836gat,G1839gat,G1840gat,G1841gat,G1844gat,G1845gat,G1846gat,G1849gat,G1850gat,G1851gat,G1854gat,G1855gat,G1856gat,G1859gat,G1860gat,G1861gat,G1864gat,G1865gat,G1866gat,G1869gat,G1870gat,G1871gat,G1874gat,G1875gat,G1876gat,G1879gat,G1880gat,G1881gat,G1884gat,G1885gat,G1886gat,G1889gat,G1890gat,G1891gat,G1894gat,G1897gat,G1902gat,G1905gat,G1908gat,G1911gat,G1914gat,G1917gat,G1920gat,G1923gat,G1926gat,G1929gat,G1932gat,G1935gat,G1938gat,G1941gat,G1945gat,G1946gat,G1947gat,G1951gat,G1955gat,G1959gat,G1963gat,G1967gat,G1971gat,G1975gat,G1979gat,G1983gat,G1987gat,G1991gat,G1995gat,G1999gat,G2000gat,G2001gat,G2004gat,G2005gat,G2006gat,G2007gat,G2008gat,G2009gat,G2010gat,G2011gat,G2012gat,G2013gat,G2014gat,G2015gat,G2016gat,G2017gat,G2018gat,G2019gat,G2020gat,G2021gat,G2022gat,G2023gat,G2024gat,G2025gat,G2026gat,G2027gat,G2028gat,G2029gat,G2030gat,G2033gat,G2037gat,G2040gat,G2043gat,G2046gat,G2049gat,G2052gat,G2055gat,G2058gat,G2061gat,G2064gat,G2067gat,G2070gat,G2073gat,G2076gat,G2080gat,G2081gat,G2082gat,G2085gat,G2089gat,G2093gat,G2097gat,G2101gat,G2105gat,G2109gat,G2113gat,G2117gat,G2121gat,G2125gat,G2129gat,G2133gat,G2137gat,G2138gat,G2139gat,G2142gat,G2145gat,G2149gat,G2150gat,G2151gat,G2154gat,G2155gat,G2156gat,G2159gat,G2160gat,G2161gat,G2164gat,G2165gat,G2166gat,G2169gat,G2170gat,G2171gat,G2174gat,G2175gat,G2176gat,G2179gat,G2180gat,G2181gat,G2184gat,G2185gat,G2186gat,G2189gat,G2190gat,G2191gat,G2194gat,G2195gat,G2196gat,G2199gat,G2200gat,G2201gat,G2204gat,G2205gat,G2206gat,G2209gat,G2210gat,G2211gat,G2214gat,G2217gat,G2221gat,G2222gat,G2224gat,G2227gat,G2230gat,G2233gat,G2236gat,G2239gat,G2242gat,G2245gat,G2248gat,G2251gat,G2254gat,G2257gat,G2260gat,G2264gat,G2265gat,G2266gat,G2269gat,G2273gat,G2277gat,G2281gat,G2285gat,G2289gat,G2293gat,G2297gat,G2301gat,G2305gat,G2309gat,G2313gat,G2317gat,G2318gat,G2319gat,G2322gat,G2326gat,G2327gat,G2328gat,G2329gat,G2330gat,G2331gat,G2332gat,G2333gat,G2334gat,G2335gat,G2336gat,G2337gat,G2338gat,G2339gat,G2340gat,G2341gat,G2342gat,G2343gat,G2344gat,G2345gat,G2346gat,G2347gat,G2348gat,G2349gat,G2350gat,G2353gat,G2357gat,G2358gat,G2359gat,G2362gat,G2365gat,G2368gat,G2371gat,G2374gat,G2377gat,G2380gat,G2383gat,G2386gat,G2389gat,G2392gat,G2395gat,G2398gat,G2402gat,G2403gat,G2404gat,G2407gat,G2410gat,G2414gat,G2418gat,G2422gat,G2426gat,G2430gat,G2434gat,G2438gat,G2442gat,G2446gat,G2450gat,G2454gat,G2458gat,G2462gat,G2463gat,G2464gat,G2467gat,G2470gat,G2474gat,G2475gat,G2476gat,G2477gat,G2478gat,G2481gat,G2482gat,G2483gat,G2486gat,G2487gat,G2488gat,G2491gat,G2492gat,G2493gat,G2496gat,G2497gat,G2498gat,G2501gat,G2502gat,G2503gat,G2506gat,G2507gat,G2508gat,G2511gat,G2512gat,G2513gat,G2516gat,G2517gat,G2518gat,G2521gat,G2522gat,G2523gat,G2526gat,G2527gat,G2528gat,G2531gat,G2532gat,G2533gat,G2536gat,G2539gat,G2543gat,G2544gat,G2545gat,G2549gat,G2552gat,G2555gat,G2558gat,G2561gat,G2564gat,G2567gat,G2570gat,G2573gat,G2576gat,G2579gat,G2582gat,G2586gat,G2587gat,G2588gat,G2591gat,G2595gat,G2599gat,G2603gat,G2607gat,G2611gat,G2615gat,G2619gat,G2623gat,G2627gat,G2631gat,G2635gat,G2639gat,G2640gat,G2641gat,G2644gat,G2648gat,G2649gat,G2650gat,G2653gat,G2654gat,G2655gat,G2656gat,G2657gat,G2658gat,G2659gat,G2660gat,G2661gat,G2662gat,G2663gat,G2664gat,G2665gat,G2666gat,G2667gat,G2668gat,G2669gat,G2670gat,G2671gat,G2672gat,G2673gat,G2674gat,G2675gat,G2678gat,G2682gat,G2683gat,G2684gat,G2687gat,G2690gat,G2694gat,G2697gat,G2700gat,G2703gat,G2706gat,G2709gat,G2712gat,G2715gat,G2718gat,G2721gat,G2724gat,G2727gat,G2731gat,G2732gat,G2733gat,G2736gat,G2739gat,G2743gat,G2744gat,G2745gat,G2749gat,G2753gat,G2757gat,G2761gat,G2765gat,G2769gat,G2773gat,G2777gat,G2781gat,G2785gat,G2789gat,G2790gat,G2791gat,G2794gat,G2797gat,G2801gat,G2802gat,G2803gat,G2806gat,G2807gat,G2808gat,G2811gat,G2812gat,G2813gat,G2816gat,G2817gat,G2818gat,G2821gat,G2822gat,G2823gat,G2826gat,G2827gat,G2828gat,G2831gat,G2832gat,G2833gat,G2836gat,G2837gat,G2838gat,G2841gat,G2842gat,G2843gat,G2846gat,G2847gat,G2848gat,G2851gat,G2852gat,G2853gat,G2856gat,G2857gat,G2858gat,G2861gat,G2864gat,G2868gat,G2869gat,G2870gat,G2873gat,G2878gat,G2881gat,G2884gat,G2887gat,G2890gat,G2893gat,G2896gat,G2899gat,G2902gat,G2905gat,G2908gat,G2912gat,G2913gat,G2914gat,G2917gat,G2921gat,G2922gat,G2923gat,G2926gat,G2930gat,G2934gat,G2938gat,G2942gat,G2946gat,G2950gat,G2954gat,G2958gat,G2962gat,G2966gat,G2967gat,G2968gat,G2971gat,G2975gat,G2976gat,G2977gat,G2980gat,G2983gat,G2987gat,G2988gat,G2989gat,G2990gat,G2991gat,G2992gat,G2993gat,G2994gat,G2995gat,G2996gat,G2997gat,G2998gat,G2999gat,G3000gat,G3001gat,G3002gat,G3003gat,G3004gat,G3005gat,G3006gat,G3007gat,G3010gat,G3014gat,G3015gat,G3016gat,G3019gat,G3022gat,G3026gat,G3027gat,G3028gat,G3031gat,G3034gat,G3037gat,G3040gat,G3043gat,G3046gat,G3049gat,G3052gat,G3055gat,G3058gat,G3062gat,G3063gat,G3064gat,G3067gat,G3070gat,G3074gat,G3075gat,G3076gat,G3079gat,G3083gat,G3087gat,G3091gat,G3095gat,G3099gat,G3103gat,G3107gat,G3111gat,G3115gat,G3119gat,G3120gat,G3121gat,G3124gat,G3127gat,G3131gat,G3132gat,G3133gat,G3136gat,G3140gat,G3141gat,G3142gat,G3145gat,G3146gat,G3147gat,G3150gat,G3151gat,G3152gat,G3155gat,G3156gat,G3157gat,G3160gat,G3161gat,G3162gat,G3165gat,G3166gat,G3167gat,G3170gat,G3171gat,G3172gat,G3175gat,G3176gat,G3177gat,G3180gat,G3181gat,G3182gat,G3185gat,G3186gat,G3187gat,G3190gat,G3193gat,G3197gat,G3198gat,G3199gat,G3202gat,G3206gat,G3207gat,G3208gat,G3212gat,G3215gat,G3218gat,G3221gat,G3224gat,G3227gat,G3230gat,G3233gat,G3236gat,G3239gat,G3243gat,G3244gat,G3245gat,G3248gat,G3252gat,G3253gat,G3254gat,G3257gat,G3260gat,G3264gat,G3268gat,G3272gat,G3276gat,G3280gat,G3284gat,G3288gat,G3292gat,G3296gat,G3300gat,G3301gat,G3302gat,G3305gat,G3309gat,G3310gat,G3311gat,G3314gat,G3317gat,G3321gat,G3322gat,G3323gat,G3324gat,G3325gat,G3326gat,G3327gat,G3328gat,G3329gat,G3330gat,G3331gat,G3332gat,G3333gat,G3334gat,G3335gat,G3336gat,G3337gat,G3338gat,G3339gat,G3340gat,G3341gat,G3344gat,G3348gat,G3349gat,G3350gat,G3353gat,G3356gat,G3360gat,G3361gat,G3362gat,G3365gat,G3368gat,G3371gat,G3374gat,G3377gat,G3380gat,G3383gat,G3386gat,G3389gat,G3392gat,G3396gat,G3397gat,G3398gat,G3401gat,G3404gat,G3408gat,G3409gat,G3410gat,G3413gat,G3417gat,G3421gat,G3425gat,G3429gat,G3433gat,G3437gat,G3441gat,G3445gat,G3449gat,G3453gat,G3454gat,G3455gat,G3458gat,G3461gat,G3465gat,G3466gat,G3467gat,G3470gat,G3474gat,G3475gat,G3476gat,G3479gat,G3480gat,G3481gat,G3484gat,G3485gat,G3486gat,G3489gat,G3490gat,G3491gat,G3494gat,G3495gat,G3496gat,G3499gat,G3500gat,G3501gat,G3504gat,G3505gat,G3506gat,G3509gat,G3510gat,G3511gat,G3514gat,G3515gat,G3516gat,G3519gat,G3520gat,G3521gat,G3524gat,G3527gat,G3531gat,G3532gat,G3533gat,G3536gat,G3540gat,G3541gat,G3542gat,G3545gat,G3548gat,G3553gat,G3556gat,G3559gat,G3562gat,G3565gat,G3568gat,G3571gat,G3574gat,G3577gat,G3581gat,G3582gat,G3583gat,G3586gat,G3590gat,G3591gat,G3592gat,G3595gat,G3598gat,G3602gat,G3603gat,G3604gat,G3608gat,G3612gat,G3616gat,G3620gat,G3624gat,G3628gat,G3632gat,G3636gat,G3637gat,G3638gat,G3641gat,G3645gat,G3646gat,G3647gat,G3650gat,G3653gat,G3657gat,G3658gat,G3659gat,G3662gat,G3663gat,G3664gat,G3665gat,G3666gat,G3667gat,G3668gat,G3669gat,G3670gat,G3671gat,G3672gat,G3673gat,G3674gat,G3675gat,G3676gat,G3677gat,G3678gat,G3681gat,G3685gat,G3686gat,G3687gat,G3690gat,G3693gat,G3697gat,G3698gat,G3699gat,G3702gat,G3706gat,G3709gat,G3712gat,G3715gat,G3718gat,G3721gat,G3724gat,G3727gat,G3730gat,G3734gat,G3735gat,G3736gat,G3739gat,G3742gat,G3746gat,G3747gat,G3748gat,G3751gat,G3755gat,G3756gat,G3757gat,G3760gat,G3764gat,G3768gat,G3772gat,G3776gat,G3780gat,G3784gat,G3788gat,G3792gat,G3793gat,G3794gat,G3797gat,G3800gat,G3804gat,G3805gat,G3806gat,G3809gat,G3813gat,G3814gat,G3815gat,G3818gat,G3821gat,G3825gat,G3826gat,G3827gat,G3830gat,G3831gat,G3832gat,G3835gat,G3836gat,G3837gat,G3840gat,G3841gat,G3842gat,G3845gat,G3846gat,G3847gat,G3850gat,G3851gat,G3852gat,G3855gat,G3856gat,G3857gat,G3860gat,G3861gat,G3862gat,G3865gat,G3868gat,G3872gat,G3873gat,G3874gat,G3877gat,G3881gat,G3882gat,G3883gat,G3886gat,G3889gat,G3893gat,G3894gat,G3896gat,G3899gat,G3902gat,G3905gat,G3908gat,G3911gat,G3914gat,G3917gat,G3921gat,G3922gat,G3923gat,G3926gat,G3930gat,G3931gat,G3932gat,G3935gat,G3938gat,G3942gat,G3943gat,G3944gat,G3947gat,G3951gat,G3955gat,G3959gat,G3963gat,G3967gat,G3971gat,G3975gat,G3976gat,G3977gat,G3980gat,G3984gat,G3985gat,G3986gat,G3989gat,G3992gat,G3996gat,G3997gat,G3998gat,G4001gat,G4005gat,G4006gat,G4007gat,G4008gat,G4009gat,G4010gat,G4011gat,G4012gat,G4013gat,G4014gat,G4015gat,G4016gat,G4017gat,G4018gat,G4019gat,G4022gat,G4026gat,G4027gat,G4028gat,G4031gat,G4034gat,G4038gat,G4039gat,G4040gat,G4043gat,G4047gat,G4048gat,G4049gat,G4052gat,G4055gat,G4058gat,G4061gat,G4064gat,G4067gat,G4070gat,G4073gat,G4077gat,G4078gat,G4079gat,G4082gat,G4085gat,G4089gat,G4090gat,G4091gat,G4094gat,G4098gat,G4099gat,G4100gat,G4103gat,G4106gat,G4110gat,G4114gat,G4118gat,G4122gat,G4126gat,G4130gat,G4134gat,G4138gat,G4139gat,G4140gat,G4143gat,G4146gat,G4150gat,G4151gat,G4152gat,G4155gat,G4159gat,G4160gat,G4161gat,G4164gat,G4167gat,G4171gat,G4172gat,G4173gat,G4174gat,G4175gat,G4178gat,G4179gat,G4180gat,G4183gat,G4184gat,G4185gat,G4188gat,G4189gat,G4190gat,G4193gat,G4194gat,G4195gat,G4198gat,G4199gat,G4200gat,G4203gat,G4204gat,G4205gat,G4208gat,G4211gat,G4215gat,G4216gat,G4217gat,G4220gat,G4224gat,G4225gat,G4226gat,G4229gat,G4232gat,G4236gat,G4237gat,G4238gat,G4242gat,G4245gat,G4248gat,G4251gat,G4254gat,G4257gat,G4260gat,G4264gat,G4265gat,G4266gat,G4269gat,G4273gat,G4274gat,G4275gat,G4278gat,G4281gat,G4285gat,G4286gat,G4287gat,G4290gat,G4294gat,G4298gat,G4302gat,G4306gat,G4310gat,G4314gat,G4318gat,G4319gat,G4320gat,G4323gat,G4327gat,G4328gat,G4329gat,G4332gat,G4335gat,G4339gat,G4340gat,G4341gat,G4344gat,G4348gat,G4349gat,G4350gat,G4353gat,G4354gat,G4355gat,G4356gat,G4357gat,G4358gat,G4359gat,G4360gat,G4361gat,G4362gat,G4363gat,G4364gat,G4365gat,G4368gat,G4372gat,G4373gat,G4374gat,G4377gat,G4380gat,G4384gat,G4385gat,G4386gat,G4389gat,G4393gat,G4394gat,G4395gat,G4398gat,G4401gat,G4405gat,G4408gat,G4411gat,G4414gat,G4417gat,G4420gat,G4423gat,G4427gat,G4428gat,G4429gat,G4432gat,G4435gat,G4439gat,G4440gat,G4441gat,G4444gat,G4448gat,G4449gat,G4450gat,G4453gat,G4456gat,G4460gat,G4461gat,G4462gat,G4466gat,G4470gat,G4474gat,G4478gat,G4482gat,G4486gat,G4487gat,G4488gat,G4491gat,G4494gat,G4498gat,G4499gat,G4500gat,G4503gat,G4507gat,G4508gat,G4509gat,G4512gat,G4515gat,G4519gat,G4520gat,G4521gat,G4524gat,G4525gat,G4526gat,G4529gat,G4530gat,G4531gat,G4534gat,G4535gat,G4536gat,G4539gat,G4540gat,G4541gat,G4544gat,G4545gat,G4546gat,G4549gat,G4550gat,G4551gat,G4554gat,G4557gat,G4561gat,G4562gat,G4563gat,G4566gat,G4570gat,G4571gat,G4572gat,G4575gat,G4578gat,G4582gat,G4583gat,G4584gat,G4587gat,G4592gat,G4595gat,G4598gat,G4601gat,G4604gat,G4607gat,G4611gat,G4612gat,G4613gat,G4616gat,G4620gat,G4621gat,G4622gat,G4625gat,G4628gat,G4632gat,G4633gat,G4634gat,G4637gat,G4641gat,G4642gat,G4643gat,G4646gat,G4650gat,G4654gat,G4658gat,G4662gat,G4666gat,G4667gat,G4668gat,G4671gat,G4675gat,G4676gat,G4677gat,G4680gat,G4683gat,G4687gat,G4688gat,G4689gat,G4692gat,G4696gat,G4697gat,G4698gat,G4701gat,G4704gat,G4708gat,G4709gat,G4710gat,G4711gat,G4712gat,G4713gat,G4714gat,G4715gat,G4716gat,G4717gat,G4718gat,G4721gat,G4725gat,G4726gat,G4727gat,G4730gat,G4733gat,G4737gat,G4738gat,G4739gat,G4742gat,G4746gat,G4747gat,G4748gat,G4751gat,G4754gat,G4758gat,G4759gat,G4760gat,G4763gat,G4766gat,G4769gat,G4772gat,G4775gat,G4779gat,G4780gat,G4781gat,G4784gat,G4787gat,G4791gat,G4792gat,G4793gat,G4796gat,G4800gat,G4801gat,G4802gat,G4805gat,G4808gat,G4812gat,G4813gat,G4814gat,G4817gat,G4821gat,G4825gat,G4829gat,G4833gat,G4837gat,G4838gat,G4839gat,G4842gat,G4845gat,G4849gat,G4850gat,G4851gat,G4854gat,G4858gat,G4859gat,G4860gat,G4863gat,G4866gat,G4870gat,G4871gat,G4872gat,G4875gat,G4879gat,G4880gat,G4881gat,G4884gat,G4885gat,G4886gat,G4889gat,G4890gat,G4891gat,G4894gat,G4895gat,G4896gat,G4899gat,G4900gat,G4901gat,G4904gat,G4907gat,G4911gat,G4912gat,G4913gat,G4916gat,G4920gat,G4921gat,G4922gat,G4925gat,G4928gat,G4932gat,G4933gat,G4934gat,G4937gat,G4941gat,G4942gat,G4943gat,G4947gat,G4950gat,G4953gat,G4956gat,G4959gat,G4963gat,G4964gat,G4965gat,G4968gat,G4972gat,G4973gat,G4974gat,G4977gat,G4980gat,G4984gat,G4985gat,G4986gat,G4989gat,G4993gat,G4994gat,G4995gat,G4998gat,G5001gat,G5005gat,G5009gat,G5013gat,G5017gat,G5021gat,G5022gat,G5023gat,G5026gat,G5030gat,G5031gat,G5032gat,G5035gat,G5038gat,G5042gat,G5043gat,G5044gat,G5047gat,G5051gat,G5052gat,G5053gat,G5056gat,G5059gat,G5063gat,G5064gat,G5065gat,G5066gat,G5067gat,G5068gat,G5069gat,G5070gat,G5071gat,G5072gat,G5073gat,G5076gat,G5080gat,G5081gat,G5082gat,G5085gat,G5088gat,G5092gat,G5093gat,G5094gat,G5097gat,G5101gat,G5102gat,G5103gat,G5106gat,G5109gat,G5113gat,G5114gat,G5115gat,G5118gat,G5121gat,G5124gat,G5127gat,G5130gat,G5134gat,G5135gat,G5136gat,G5139gat,G5142gat,G5146gat,G5147gat,G5148gat,G5151gat,G5155gat,G5156gat,G5157gat,G5160gat,G5163gat,G5167gat,G5168gat,G5169gat,G5172gat,G5176gat,G5180gat,G5184gat,G5188gat,G5192gat,G5193gat,G5194gat,G5197gat,G5200gat,G5204gat,G5205gat,G5206gat,G5209gat,G5213gat,G5214gat,G5215gat,G5218gat,G5221gat,G5225gat,G5226gat,G5227gat,G5230gat,G5234gat,G5235gat,G5236gat,G5239gat,G5240gat,G5241gat,G5244gat,G5245gat,G5246gat,G5249gat,G5250gat,G5251gat,G5254gat,G5255gat,G5256gat,G5259gat,G5262gat,G5266gat,G5267gat,G5268gat,G5271gat,G5275gat,G5276gat,G5277gat,G5280gat,G5283gat,G5287gat,G5288gat,G5289gat,G5292gat,G5296gat,G5297gat,G5298gat,G5301gat,G5304gat,G5309gat,G5312gat,G5315gat,G5318gat,G5322gat,G5323gat,G5324gat,G5327gat,G5331gat,G5332gat,G5333gat,G5336gat,G5339gat,G5343gat,G5344gat,G5345gat,G5348gat,G5352gat,G5353gat,G5354gat,G5357gat,G5360gat,G5364gat,G5365gat,G5366gat,G5370gat,G5374gat,G5378gat,G5379gat,G5380gat,G5383gat,G5387gat,G5388gat,G5389gat,G5392gat,G5395gat,G5399gat,G5400gat,G5401gat,G5404gat,G5408gat,G5409gat,G5410gat,G5413gat,G5416gat,G5420gat,G5421gat,G5422gat,G5425gat,G5426gat,G5427gat,G5428gat,G5429gat,G5430gat,G5431gat,G5434gat,G5438gat,G5439gat,G5440gat,G5443gat,G5446gat,G5450gat,G5451gat,G5452gat,G5455gat,G5459gat,G5460gat,G5461gat,G5464gat,G5467gat,G5471gat,G5472gat,G5473gat,G5476gat,G5480gat,G5483gat,G5486gat,G5489gat,G5493gat,G5494gat,G5495gat,G5498gat,G5501gat,G5505gat,G5506gat,G5507gat,G5510gat,G5514gat,G5515gat,G5516gat,G5519gat,G5522gat,G5526gat,G5527gat,G5528gat,G5531gat,G5535gat,G5536gat,G5537gat,G5540gat,G5544gat,G5548gat,G5552gat,G5553gat,G5554gat,G5557gat,G5560gat,G5564gat,G5565gat,G5566gat,G5569gat,G5573gat,G5574gat,G5575gat,G5578gat,G5581gat,G5585gat,G5586gat,G5587gat,G5590gat,G5594gat,G5595gat,G5596gat,G5599gat,G5602gat,G5606gat,G5607gat,G5608gat,G5611gat,G5612gat,G5613gat,G5616gat,G5617gat,G5618gat,G5621gat,G5624gat,G5628gat,G5629gat,G5630gat,G5633gat,G5637gat,G5638gat,G5639gat,G5642gat,G5645gat,G5649gat,G5650gat,G5651gat,G5654gat,G5658gat,G5659gat,G5660gat,G5663gat,G5666gat,G5670gat,G5671gat,G5673gat,G5676gat,G5679gat,G5683gat,G5684gat,G5685gat,G5688gat,G5692gat,G5693gat,G5694gat,G5697gat,G5700gat,G5704gat,G5705gat,G5706gat,G5709gat,G5713gat,G5714gat,G5715gat,G5718gat,G5721gat,G5725gat,G5726gat,G5727gat,G5730gat,G5734gat,G5738gat,G5739gat,G5740gat,G5743gat,G5747gat,G5748gat,G5749gat,G5752gat,G5755gat,G5759gat,G5760gat,G5761gat,G5764gat,G5768gat,G5769gat,G5770gat,G5773gat,G5776gat,G5780gat,G5781gat,G5782gat,G5785gat,G5786gat,G5787gat,G5788gat,G5789gat,G5792gat,G5796gat,G5797gat,G5798gat,G5801gat,G5804gat,G5808gat,G5809gat,G5810gat,G5813gat,G5817gat,G5818gat,G5819gat,G5822gat,G5825gat,G5829gat,G5830gat,G5831gat,G5834gat,G5837gat,G5840gat,G5844gat,G5845gat,G5846gat,G5849gat,G5852gat,G5856gat,G5857gat,G5858gat,G5861gat,G5865gat,G5866gat,G5867gat,G5870gat,G5873gat,G5877gat,G5878gat,G5879gat,G5882gat,G5886gat,G5890gat,G5891gat,G5892gat,G5895gat,G5898gat,G5902gat,G5903gat,G5904gat,G5907gat,G5911gat,G5912gat,G5913gat,G5916gat,G5919gat,G5923gat,G5924gat,G5925gat,G5928gat,G5929gat,G5930gat,G5933gat,G5934gat,G5935gat,G5938gat,G5941gat,G5945gat,G5946gat,G5947gat,G5950gat,G5954gat,G5955gat,G5956gat,G5959gat,G5962gat,G5966gat,G5967gat,G5968gat,G5972gat,G5975gat,G5979gat,G5980gat,G5981gat,G5984gat,G5988gat,G5989gat,G5990gat,G5993gat,G5996gat,G6000gat,G6001gat,G6002gat,G6005gat,G6009gat,G6010gat,G6011gat,G6014gat,G6018gat,G6019gat,G6020gat,G6023gat,G6026gat,G6030gat,G6031gat,G6032gat,G6035gat,G6036gat,G6037gat,G6040gat,G6044gat,G6045gat,G6046gat,G6049gat,G6052gat,G6056gat,G6057gat,G6058gat,G6061gat,G6064gat,G6068gat,G6069gat,G6070gat,G6073gat,G6076gat,G6080gat,G6081gat,G6082gat,G6085gat,G6089gat,G6090gat,G6091gat,G6094gat,G6097gat,G6101gat,G6102gat,G6103gat,G6106gat,G6107gat,G6108gat,G6111gat,G6114gat,G6118gat,G6119gat,G6120gat,G6124gat,G6128gat,G6129gat,G6130gat,G6133gat,G6134gat,G6135gat,G6138gat,G6141gat,G6145gat,G6146gat,G6147gat,G6151gat,G6155gat,G6156gat,G6157gat,G6161gat,G6165gat,G6166gat,G6167gat,G6171gat,G6175gat,G6176gat,G6177gat,G6181gat,G6185gat,G6186gat,G6187gat,G6191gat,G6195gat,G6196gat,G6197gat,G6201gat,G6205gat,G6206gat,G6207gat,G6211gat,G6215gat,G6216gat,G6217gat,G6221gat,G6225gat,G6226gat,G6227gat,G6231gat,G6235gat,G6236gat,G6237gat,G6241gat,G6245gat,G6246gat,G6247gat,G6251gat,G6255gat,G6256gat,G6257gat,G6261gat,G6265gat,G6266gat,G6267gat,G6271gat,G6275gat,G6276gat,G6277gat,G6281gat,G6285gat,G6286gat;

and AND2_1 (G545gat, G1gat, G273gat);
and AND2_2 (G546gat, G1gat, G290gat);
and AND2_3 (G549gat_enc, G1gat, G307gat);
xnor XNOR2_4 (G549gat, keyinput0, G549gat_enc);
and AND2_5 (G552gat, G1gat, G324gat);
and AND2_6 (G555gat_enc, G1gat, G341gat);
xnor XNOR2_7 (G555gat, keyinput1, G555gat_enc);
and AND2_8 (G558gat_enc, G1gat, G358gat);
nor NOR2_9 (CLK8, G558gat_enc, G555gat);
dff DFF2_10 (LIBAR8, CLK8, keyinput2);
xor XOR2_11 (G558gat, LIBAR8, G558gat_enc);
and AND2_12 (G561gat_enc, G1gat, G375gat);
xor XOR2_13 (G561gat, keyinput3, G561gat_enc);
and AND2_14 (G564gat_enc, G1gat, G392gat);
xor XOR2_15 (G564gat, keyinput4, G564gat_enc);
and AND2_16 (G567gat, G1gat, G409gat);
and AND2_17 (G570gat_enc, G1gat, G426gat);
xnor XNOR2_18 (G570gat, keyinput5, G570gat_enc);
and AND2_19 (G573gat_enc, G1gat, G443gat);
xnor XNOR2_20 (G573gat, keyinput6, G573gat_enc);
and AND2_21 (G576gat_enc, G1gat, G460gat);
xor XOR2_22 (G576gat, keyinput7, G576gat_enc);
and AND2_23 (G579gat_enc, G1gat, G477gat);
nor NOR2_24 (CLK7, G579gat_enc, G576gat);
dff DFF2_25 (LIBAR7, CLK7, keyinput8);
xnor XNOR2_26 (G579gat, LIBAR7, G579gat_enc);
and AND2_27 (G582gat_enc, G1gat, G494gat);
xor XOR2_28 (G582gat, keyinput9, G582gat_enc);
and AND2_29 (G585gat, G1gat, G511gat);
and AND2_30 (G588gat, G1gat, G528gat);
and AND2_31 (G591gat_enc, G18gat, G273gat);
nor NOR2_32 (CLK6, G591gat_enc, G588gat);
dff DFF2_33 (LIBAR6, CLK6, keyinput10);
xnor XNOR2_34 (G591gat, LIBAR6, G591gat_enc);
and AND2_35 (G594gat_enc, G18gat, G290gat);
nor NOR2_36 (CLK5, G594gat_enc, G591gat);
dff DFF2_37 (LIBAR5, CLK5, keyinput11);
xor XOR2_38 (G594gat, LIBAR5, G594gat_enc);
and AND2_39 (G597gat_enc, G18gat, G307gat);
nor NOR2_40 (CLK4, G597gat_enc, G594gat);
dff DFF2_41 (LIBAR4, CLK4, keyinput12);
xnor XNOR2_42 (G597gat, LIBAR4, G597gat_enc);
and AND2_43 (G600gat, G18gat, G324gat);
and AND2_44 (G603gat, G18gat, G341gat);
and AND2_45 (G606gat_enc, G18gat, G358gat);
nor NOR2_46 (CLK3, G606gat_enc, G603gat);
dff DFF2_47 (LIBAR3, CLK3, keyinput13);
xnor XNOR2_48 (G606gat, LIBAR3, G606gat_enc);
and AND2_49 (G609gat_enc, G18gat, G375gat);
nor NOR2_50 (CLK2, G609gat_enc, G606gat);
dff DFF2_51 (LIBAR2, CLK2, keyinput14);
xor XOR2_52 (G609gat, LIBAR2, G609gat_enc);
and AND2_53 (G612gat_enc, G18gat, G392gat);
nor NOR2_54 (CLK1, G612gat_enc, G609gat);
dff DFF2_55 (LIBAR1, CLK1, keyinput15);
xor XOR2_56 (G612gat, LIBAR1, G612gat_enc);
and AND2_57 (G615gat, G18gat, G409gat);
and AND2_58 (G618gat, G18gat, G426gat);
and AND2_59 (G621gat, G18gat, G443gat);
and AND2_60 (G624gat, G18gat, G460gat);
and AND2_61 (G627gat, G18gat, G477gat);
and AND2_62 (G630gat, G18gat, G494gat);
and AND2_63 (G633gat, G18gat, G511gat);
and AND2_64 (G636gat, G18gat, G528gat);
and AND2_65 (G639gat, G35gat, G273gat);
and AND2_66 (G642gat, G35gat, G290gat);
and AND2_67 (G645gat, G35gat, G307gat);
and AND2_68 (G648gat, G35gat, G324gat);
and AND2_69 (G651gat, G35gat, G341gat);
and AND2_70 (G654gat, G35gat, G358gat);
and AND2_71 (G657gat, G35gat, G375gat);
and AND2_72 (G660gat, G35gat, G392gat);
and AND2_73 (G663gat, G35gat, G409gat);
and AND2_74 (G666gat, G35gat, G426gat);
and AND2_75 (G669gat, G35gat, G443gat);
and AND2_76 (G672gat, G35gat, G460gat);
and AND2_77 (G675gat, G35gat, G477gat);
and AND2_78 (G678gat, G35gat, G494gat);
and AND2_79 (G681gat, G35gat, G511gat);
and AND2_80 (G684gat, G35gat, G528gat);
and AND2_81 (G687gat, G52gat, G273gat);
and AND2_82 (G690gat, G52gat, G290gat);
and AND2_83 (G693gat, G52gat, G307gat);
and AND2_84 (G696gat, G52gat, G324gat);
and AND2_85 (G699gat, G52gat, G341gat);
and AND2_86 (G702gat, G52gat, G358gat);
and AND2_87 (G705gat, G52gat, G375gat);
and AND2_88 (G708gat, G52gat, G392gat);
and AND2_89 (G711gat, G52gat, G409gat);
and AND2_90 (G714gat, G52gat, G426gat);
and AND2_91 (G717gat, G52gat, G443gat);
and AND2_92 (G720gat, G52gat, G460gat);
and AND2_93 (G723gat, G52gat, G477gat);
and AND2_94 (G726gat, G52gat, G494gat);
and AND2_95 (G729gat, G52gat, G511gat);
and AND2_96 (G732gat, G52gat, G528gat);
and AND2_97 (G735gat, G69gat, G273gat);
and AND2_98 (G738gat, G69gat, G290gat);
and AND2_99 (G741gat, G69gat, G307gat);
and AND2_100 (G744gat, G69gat, G324gat);
and AND2_101 (G747gat, G69gat, G341gat);
and AND2_102 (G750gat, G69gat, G358gat);
and AND2_103 (G753gat, G69gat, G375gat);
and AND2_104 (G756gat, G69gat, G392gat);
and AND2_105 (G759gat, G69gat, G409gat);
and AND2_106 (G762gat, G69gat, G426gat);
and AND2_107 (G765gat, G69gat, G443gat);
and AND2_108 (G768gat, G69gat, G460gat);
and AND2_109 (G771gat, G69gat, G477gat);
and AND2_110 (G774gat, G69gat, G494gat);
and AND2_111 (G777gat, G69gat, G511gat);
and AND2_112 (G780gat, G69gat, G528gat);
and AND2_113 (G783gat, G86gat, G273gat);
and AND2_114 (G786gat, G86gat, G290gat);
and AND2_115 (G789gat, G86gat, G307gat);
and AND2_116 (G792gat, G86gat, G324gat);
and AND2_117 (G795gat, G86gat, G341gat);
and AND2_118 (G798gat, G86gat, G358gat);
and AND2_119 (G801gat, G86gat, G375gat);
and AND2_120 (G804gat, G86gat, G392gat);
and AND2_121 (G807gat, G86gat, G409gat);
and AND2_122 (G810gat, G86gat, G426gat);
and AND2_123 (G813gat, G86gat, G443gat);
and AND2_124 (G816gat, G86gat, G460gat);
and AND2_125 (G819gat, G86gat, G477gat);
and AND2_126 (G822gat, G86gat, G494gat);
and AND2_127 (G825gat, G86gat, G511gat);
and AND2_128 (G828gat, G86gat, G528gat);
and AND2_129 (G831gat, G103gat, G273gat);
and AND2_130 (G834gat, G103gat, G290gat);
and AND2_131 (G837gat, G103gat, G307gat);
and AND2_132 (G840gat, G103gat, G324gat);
and AND2_133 (G843gat, G103gat, G341gat);
and AND2_134 (G846gat, G103gat, G358gat);
and AND2_135 (G849gat, G103gat, G375gat);
and AND2_136 (G852gat, G103gat, G392gat);
and AND2_137 (G855gat, G103gat, G409gat);
and AND2_138 (G858gat, G103gat, G426gat);
and AND2_139 (G861gat, G103gat, G443gat);
and AND2_140 (G864gat, G103gat, G460gat);
and AND2_141 (G867gat, G103gat, G477gat);
and AND2_142 (G870gat, G103gat, G494gat);
and AND2_143 (G873gat, G103gat, G511gat);
and AND2_144 (G876gat, G103gat, G528gat);
and AND2_145 (G879gat, G120gat, G273gat);
and AND2_146 (G882gat, G120gat, G290gat);
and AND2_147 (G885gat, G120gat, G307gat);
and AND2_148 (G888gat, G120gat, G324gat);
and AND2_149 (G891gat, G120gat, G341gat);
and AND2_150 (G894gat, G120gat, G358gat);
and AND2_151 (G897gat, G120gat, G375gat);
and AND2_152 (G900gat, G120gat, G392gat);
and AND2_153 (G903gat, G120gat, G409gat);
and AND2_154 (G906gat, G120gat, G426gat);
and AND2_155 (G909gat, G120gat, G443gat);
and AND2_156 (G912gat, G120gat, G460gat);
and AND2_157 (G915gat, G120gat, G477gat);
and AND2_158 (G918gat, G120gat, G494gat);
and AND2_159 (G921gat, G120gat, G511gat);
and AND2_160 (G924gat, G120gat, G528gat);
and AND2_161 (G927gat, G137gat, G273gat);
and AND2_162 (G930gat, G137gat, G290gat);
and AND2_163 (G933gat, G137gat, G307gat);
and AND2_164 (G936gat, G137gat, G324gat);
and AND2_165 (G939gat, G137gat, G341gat);
and AND2_166 (G942gat, G137gat, G358gat);
and AND2_167 (G945gat, G137gat, G375gat);
and AND2_168 (G948gat, G137gat, G392gat);
and AND2_169 (G951gat, G137gat, G409gat);
and AND2_170 (G954gat, G137gat, G426gat);
and AND2_171 (G957gat, G137gat, G443gat);
and AND2_172 (G960gat, G137gat, G460gat);
and AND2_173 (G963gat, G137gat, G477gat);
and AND2_174 (G966gat, G137gat, G494gat);
and AND2_175 (G969gat, G137gat, G511gat);
and AND2_176 (G972gat, G137gat, G528gat);
and AND2_177 (G975gat, G154gat, G273gat);
and AND2_178 (G978gat, G154gat, G290gat);
and AND2_179 (G981gat, G154gat, G307gat);
and AND2_180 (G984gat, G154gat, G324gat);
and AND2_181 (G987gat, G154gat, G341gat);
and AND2_182 (G990gat, G154gat, G358gat);
and AND2_183 (G993gat, G154gat, G375gat);
and AND2_184 (G996gat, G154gat, G392gat);
and AND2_185 (G999gat, G154gat, G409gat);
and AND2_186 (G1002gat, G154gat, G426gat);
and AND2_187 (G1005gat, G154gat, G443gat);
and AND2_188 (G1008gat, G154gat, G460gat);
and AND2_189 (G1011gat, G154gat, G477gat);
and AND2_190 (G1014gat, G154gat, G494gat);
and AND2_191 (G1017gat, G154gat, G511gat);
and AND2_192 (G1020gat, G154gat, G528gat);
and AND2_193 (G1023gat, G171gat, G273gat);
and AND2_194 (G1026gat, G171gat, G290gat);
and AND2_195 (G1029gat, G171gat, G307gat);
and AND2_196 (G1032gat, G171gat, G324gat);
and AND2_197 (G1035gat, G171gat, G341gat);
and AND2_198 (G1038gat, G171gat, G358gat);
and AND2_199 (G1041gat, G171gat, G375gat);
and AND2_200 (G1044gat, G171gat, G392gat);
and AND2_201 (G1047gat, G171gat, G409gat);
and AND2_202 (G1050gat, G171gat, G426gat);
and AND2_203 (G1053gat, G171gat, G443gat);
and AND2_204 (G1056gat, G171gat, G460gat);
and AND2_205 (G1059gat, G171gat, G477gat);
and AND2_206 (G1062gat, G171gat, G494gat);
and AND2_207 (G1065gat, G171gat, G511gat);
and AND2_208 (G1068gat, G171gat, G528gat);
and AND2_209 (G1071gat, G188gat, G273gat);
and AND2_210 (G1074gat, G188gat, G290gat);
and AND2_211 (G1077gat, G188gat, G307gat);
and AND2_212 (G1080gat, G188gat, G324gat);
and AND2_213 (G1083gat, G188gat, G341gat);
and AND2_214 (G1086gat, G188gat, G358gat);
and AND2_215 (G1089gat, G188gat, G375gat);
and AND2_216 (G1092gat, G188gat, G392gat);
and AND2_217 (G1095gat, G188gat, G409gat);
and AND2_218 (G1098gat, G188gat, G426gat);
and AND2_219 (G1101gat, G188gat, G443gat);
and AND2_220 (G1104gat, G188gat, G460gat);
and AND2_221 (G1107gat, G188gat, G477gat);
and AND2_222 (G1110gat, G188gat, G494gat);
and AND2_223 (G1113gat, G188gat, G511gat);
and AND2_224 (G1116gat, G188gat, G528gat);
and AND2_225 (G1119gat, G205gat, G273gat);
and AND2_226 (G1122gat, G205gat, G290gat);
and AND2_227 (G1125gat, G205gat, G307gat);
and AND2_228 (G1128gat, G205gat, G324gat);
and AND2_229 (G1131gat, G205gat, G341gat);
and AND2_230 (G1134gat, G205gat, G358gat);
and AND2_231 (G1137gat, G205gat, G375gat);
and AND2_232 (G1140gat, G205gat, G392gat);
and AND2_233 (G1143gat, G205gat, G409gat);
and AND2_234 (G1146gat, G205gat, G426gat);
and AND2_235 (G1149gat, G205gat, G443gat);
and AND2_236 (G1152gat, G205gat, G460gat);
and AND2_237 (G1155gat, G205gat, G477gat);
and AND2_238 (G1158gat, G205gat, G494gat);
and AND2_239 (G1161gat, G205gat, G511gat);
and AND2_240 (G1164gat, G205gat, G528gat);
and AND2_241 (G1167gat, G222gat, G273gat);
and AND2_242 (G1170gat, G222gat, G290gat);
and AND2_243 (G1173gat, G222gat, G307gat);
and AND2_244 (G1176gat, G222gat, G324gat);
and AND2_245 (G1179gat, G222gat, G341gat);
and AND2_246 (G1182gat, G222gat, G358gat);
and AND2_247 (G1185gat, G222gat, G375gat);
and AND2_248 (G1188gat, G222gat, G392gat);
and AND2_249 (G1191gat, G222gat, G409gat);
and AND2_250 (G1194gat, G222gat, G426gat);
and AND2_251 (G1197gat, G222gat, G443gat);
and AND2_252 (G1200gat, G222gat, G460gat);
and AND2_253 (G1203gat, G222gat, G477gat);
and AND2_254 (G1206gat, G222gat, G494gat);
and AND2_255 (G1209gat, G222gat, G511gat);
and AND2_256 (G1212gat, G222gat, G528gat);
and AND2_257 (G1215gat, G239gat, G273gat);
and AND2_258 (G1218gat, G239gat, G290gat);
and AND2_259 (G1221gat, G239gat, G307gat);
and AND2_260 (G1224gat, G239gat, G324gat);
and AND2_261 (G1227gat, G239gat, G341gat);
and AND2_262 (G1230gat, G239gat, G358gat);
and AND2_263 (G1233gat, G239gat, G375gat);
and AND2_264 (G1236gat, G239gat, G392gat);
and AND2_265 (G1239gat, G239gat, G409gat);
and AND2_266 (G1242gat, G239gat, G426gat);
and AND2_267 (G1245gat, G239gat, G443gat);
and AND2_268 (G1248gat, G239gat, G460gat);
and AND2_269 (G1251gat, G239gat, G477gat);
and AND2_270 (G1254gat, G239gat, G494gat);
and AND2_271 (G1257gat, G239gat, G511gat);
and AND2_272 (G1260gat, G239gat, G528gat);
and AND2_273 (G1263gat, G256gat, G273gat);
and AND2_274 (G1266gat, G256gat, G290gat);
and AND2_275 (G1269gat, G256gat, G307gat);
and AND2_276 (G1272gat, G256gat, G324gat);
and AND2_277 (G1275gat, G256gat, G341gat);
and AND2_278 (G1278gat, G256gat, G358gat);
and AND2_279 (G1281gat, G256gat, G375gat);
and AND2_280 (G1284gat, G256gat, G392gat);
and AND2_281 (G1287gat, G256gat, G409gat);
and AND2_282 (G1290gat, G256gat, G426gat);
and AND2_283 (G1293gat, G256gat, G443gat);
and AND2_284 (G1296gat, G256gat, G460gat);
and AND2_285 (G1299gat, G256gat, G477gat);
and AND2_286 (G1302gat, G256gat, G494gat);
and AND2_287 (G1305gat, G256gat, G511gat);
and AND2_288 (G1308gat, G256gat, G528gat);
not NOT1_289 (G1311gat, G591gat);
not NOT1_290 (G1315gat, G639gat);
not NOT1_291 (G1319gat, G687gat);
not NOT1_292 (G1323gat, G735gat);
not NOT1_293 (G1327gat, G783gat);
not NOT1_294 (G1331gat, G831gat);
not NOT1_295 (G1335gat, G879gat);
not NOT1_296 (G1339gat, G927gat);
not NOT1_297 (G1343gat, G975gat);
not NOT1_298 (G1347gat, G1023gat);
not NOT1_299 (G1351gat, G1071gat);
not NOT1_300 (G1355gat, G1119gat);
not NOT1_301 (G1359gat, G1167gat);
not NOT1_302 (G1363gat, G1215gat);
not NOT1_303 (G1367gat, G1263gat);
nor NOR2_304 (G1371gat, G591gat, G1311gat);
not NOT1_305 (G1372gat, G1311gat);
nor NOR2_306 (G1373gat, G639gat, G1315gat);
not NOT1_307 (G1374gat, G1315gat);
nor NOR2_308 (G1375gat, G687gat, G1319gat);
not NOT1_309 (G1376gat, G1319gat);
nor NOR2_310 (G1377gat, G735gat, G1323gat);
not NOT1_311 (G1378gat, G1323gat);
nor NOR2_312 (G1379gat, G783gat, G1327gat);
not NOT1_313 (G1380gat, G1327gat);
nor NOR2_314 (G1381gat, G831gat, G1331gat);
not NOT1_315 (G1382gat, G1331gat);
nor NOR2_316 (G1383gat, G879gat, G1335gat);
not NOT1_317 (G1384gat, G1335gat);
nor NOR2_318 (G1385gat, G927gat, G1339gat);
not NOT1_319 (G1386gat, G1339gat);
nor NOR2_320 (G1387gat, G975gat, G1343gat);
not NOT1_321 (G1388gat, G1343gat);
nor NOR2_322 (G1389gat, G1023gat, G1347gat);
not NOT1_323 (G1390gat, G1347gat);
nor NOR2_324 (G1391gat, G1071gat, G1351gat);
not NOT1_325 (G1392gat, G1351gat);
nor NOR2_326 (G1393gat, G1119gat, G1355gat);
not NOT1_327 (G1394gat, G1355gat);
nor NOR2_328 (G1395gat, G1167gat, G1359gat);
not NOT1_329 (G1396gat, G1359gat);
nor NOR2_330 (G1397gat, G1215gat, G1363gat);
not NOT1_331 (G1398gat, G1363gat);
nor NOR2_332 (G1399gat, G1263gat, G1367gat);
not NOT1_333 (G1400gat, G1367gat);
nor NOR2_334 (G1401gat, G1371gat, G1372gat);
nor NOR2_335 (G1404gat, G1373gat, G1374gat);
nor NOR2_336 (G1407gat, G1375gat, G1376gat);
nor NOR2_337 (G1410gat, G1377gat, G1378gat);
nor NOR2_338 (G1413gat, G1379gat, G1380gat);
nor NOR2_339 (G1416gat, G1381gat, G1382gat);
nor NOR2_340 (G1419gat, G1383gat, G1384gat);
nor NOR2_341 (G1422gat, G1385gat, G1386gat);
nor NOR2_342 (G1425gat, G1387gat, G1388gat);
nor NOR2_343 (G1428gat, G1389gat, G1390gat);
nor NOR2_344 (G1431gat, G1391gat, G1392gat);
nor NOR2_345 (G1434gat, G1393gat, G1394gat);
nor NOR2_346 (G1437gat, G1395gat, G1396gat);
nor NOR2_347 (G1440gat, G1397gat, G1398gat);
nor NOR2_348 (G1443gat, G1399gat, G1400gat);
nor NOR2_349 (G1446gat, G1401gat, G546gat);
nor NOR2_350 (G1450gat, G1404gat, G594gat);
nor NOR2_351 (G1454gat, G1407gat, G642gat);
nor NOR2_352 (G1458gat, G1410gat, G690gat);
nor NOR2_353 (G1462gat, G1413gat, G738gat);
nor NOR2_354 (G1466gat, G1416gat, G786gat);
nor NOR2_355 (G1470gat, G1419gat, G834gat);
nor NOR2_356 (G1474gat, G1422gat, G882gat);
nor NOR2_357 (G1478gat, G1425gat, G930gat);
nor NOR2_358 (G1482gat, G1428gat, G978gat);
nor NOR2_359 (G1486gat, G1431gat, G1026gat);
nor NOR2_360 (G1490gat, G1434gat, G1074gat);
nor NOR2_361 (G1494gat, G1437gat, G1122gat);
nor NOR2_362 (G1498gat, G1440gat, G1170gat);
nor NOR2_363 (G1502gat, G1443gat, G1218gat);
nor NOR2_364 (G1506gat, G1401gat, G1446gat);
nor NOR2_365 (G1507gat, G1446gat, G546gat);
nor NOR2_366 (G1508gat, G1311gat, G1446gat);
nor NOR2_367 (G1511gat, G1404gat, G1450gat);
nor NOR2_368 (G1512gat, G1450gat, G594gat);
nor NOR2_369 (G1513gat, G1315gat, G1450gat);
nor NOR2_370 (G1516gat, G1407gat, G1454gat);
nor NOR2_371 (G1517gat, G1454gat, G642gat);
nor NOR2_372 (G1518gat, G1319gat, G1454gat);
nor NOR2_373 (G1521gat, G1410gat, G1458gat);
nor NOR2_374 (G1522gat, G1458gat, G690gat);
nor NOR2_375 (G1523gat, G1323gat, G1458gat);
nor NOR2_376 (G1526gat, G1413gat, G1462gat);
nor NOR2_377 (G1527gat, G1462gat, G738gat);
nor NOR2_378 (G1528gat, G1327gat, G1462gat);
nor NOR2_379 (G1531gat, G1416gat, G1466gat);
nor NOR2_380 (G1532gat, G1466gat, G786gat);
nor NOR2_381 (G1533gat, G1331gat, G1466gat);
nor NOR2_382 (G1536gat, G1419gat, G1470gat);
nor NOR2_383 (G1537gat, G1470gat, G834gat);
nor NOR2_384 (G1538gat, G1335gat, G1470gat);
nor NOR2_385 (G1541gat, G1422gat, G1474gat);
nor NOR2_386 (G1542gat, G1474gat, G882gat);
nor NOR2_387 (G1543gat, G1339gat, G1474gat);
nor NOR2_388 (G1546gat, G1425gat, G1478gat);
nor NOR2_389 (G1547gat, G1478gat, G930gat);
nor NOR2_390 (G1548gat, G1343gat, G1478gat);
nor NOR2_391 (G1551gat, G1428gat, G1482gat);
nor NOR2_392 (G1552gat, G1482gat, G978gat);
nor NOR2_393 (G1553gat, G1347gat, G1482gat);
nor NOR2_394 (G1556gat, G1431gat, G1486gat);
nor NOR2_395 (G1557gat, G1486gat, G1026gat);
nor NOR2_396 (G1558gat, G1351gat, G1486gat);
nor NOR2_397 (G1561gat, G1434gat, G1490gat);
nor NOR2_398 (G1562gat, G1490gat, G1074gat);
nor NOR2_399 (G1563gat, G1355gat, G1490gat);
nor NOR2_400 (G1566gat, G1437gat, G1494gat);
nor NOR2_401 (G1567gat, G1494gat, G1122gat);
nor NOR2_402 (G1568gat, G1359gat, G1494gat);
nor NOR2_403 (G1571gat, G1440gat, G1498gat);
nor NOR2_404 (G1572gat, G1498gat, G1170gat);
nor NOR2_405 (G1573gat, G1363gat, G1498gat);
nor NOR2_406 (G1576gat, G1443gat, G1502gat);
nor NOR2_407 (G1577gat, G1502gat, G1218gat);
nor NOR2_408 (G1578gat, G1367gat, G1502gat);
nor NOR2_409 (G1581gat, G1506gat, G1507gat);
nor NOR2_410 (G1582gat, G1511gat, G1512gat);
nor NOR2_411 (G1585gat, G1516gat, G1517gat);
nor NOR2_412 (G1588gat, G1521gat, G1522gat);
nor NOR2_413 (G1591gat, G1526gat, G1527gat);
nor NOR2_414 (G1594gat, G1531gat, G1532gat);
nor NOR2_415 (G1597gat, G1536gat, G1537gat);
nor NOR2_416 (G1600gat, G1541gat, G1542gat);
nor NOR2_417 (G1603gat, G1546gat, G1547gat);
nor NOR2_418 (G1606gat, G1551gat, G1552gat);
nor NOR2_419 (G1609gat, G1556gat, G1557gat);
nor NOR2_420 (G1612gat, G1561gat, G1562gat);
nor NOR2_421 (G1615gat, G1566gat, G1567gat);
nor NOR2_422 (G1618gat, G1571gat, G1572gat);
nor NOR2_423 (G1621gat, G1576gat, G1577gat);
nor NOR2_424 (G1624gat, G1266gat, G1578gat);
nor NOR2_425 (G1628gat, G1582gat, G1508gat);
nor NOR2_426 (G1632gat, G1585gat, G1513gat);
nor NOR2_427 (G1636gat, G1588gat, G1518gat);
nor NOR2_428 (G1640gat, G1591gat, G1523gat);
nor NOR2_429 (G1644gat, G1594gat, G1528gat);
nor NOR2_430 (G1648gat, G1597gat, G1533gat);
nor NOR2_431 (G1652gat, G1600gat, G1538gat);
nor NOR2_432 (G1656gat, G1603gat, G1543gat);
nor NOR2_433 (G1660gat, G1606gat, G1548gat);
nor NOR2_434 (G1664gat, G1609gat, G1553gat);
nor NOR2_435 (G1668gat, G1612gat, G1558gat);
nor NOR2_436 (G1672gat, G1615gat, G1563gat);
nor NOR2_437 (G1676gat, G1618gat, G1568gat);
nor NOR2_438 (G1680gat, G1621gat, G1573gat);
nor NOR2_439 (G1684gat, G1266gat, G1624gat);
nor NOR2_440 (G1685gat, G1624gat, G1578gat);
nor NOR2_441 (G1686gat, G1582gat, G1628gat);
nor NOR2_442 (G1687gat, G1628gat, G1508gat);
nor NOR2_443 (G1688gat, G1585gat, G1632gat);
nor NOR2_444 (G1689gat, G1632gat, G1513gat);
nor NOR2_445 (G1690gat, G1588gat, G1636gat);
nor NOR2_446 (G1691gat, G1636gat, G1518gat);
nor NOR2_447 (G1692gat, G1591gat, G1640gat);
nor NOR2_448 (G1693gat, G1640gat, G1523gat);
nor NOR2_449 (G1694gat, G1594gat, G1644gat);
nor NOR2_450 (G1695gat, G1644gat, G1528gat);
nor NOR2_451 (G1696gat, G1597gat, G1648gat);
nor NOR2_452 (G1697gat, G1648gat, G1533gat);
nor NOR2_453 (G1698gat, G1600gat, G1652gat);
nor NOR2_454 (G1699gat, G1652gat, G1538gat);
nor NOR2_455 (G1700gat, G1603gat, G1656gat);
nor NOR2_456 (G1701gat, G1656gat, G1543gat);
nor NOR2_457 (G1702gat, G1606gat, G1660gat);
nor NOR2_458 (G1703gat, G1660gat, G1548gat);
nor NOR2_459 (G1704gat, G1609gat, G1664gat);
nor NOR2_460 (G1705gat, G1664gat, G1553gat);
nor NOR2_461 (G1706gat, G1612gat, G1668gat);
nor NOR2_462 (G1707gat, G1668gat, G1558gat);
nor NOR2_463 (G1708gat, G1615gat, G1672gat);
nor NOR2_464 (G1709gat, G1672gat, G1563gat);
nor NOR2_465 (G1710gat, G1618gat, G1676gat);
nor NOR2_466 (G1711gat, G1676gat, G1568gat);
nor NOR2_467 (G1712gat, G1621gat, G1680gat);
nor NOR2_468 (G1713gat, G1680gat, G1573gat);
nor NOR2_469 (G1714gat, G1684gat, G1685gat);
nor NOR2_470 (G1717gat, G1686gat, G1687gat);
nor NOR2_471 (G1720gat, G1688gat, G1689gat);
nor NOR2_472 (G1723gat, G1690gat, G1691gat);
nor NOR2_473 (G1726gat, G1692gat, G1693gat);
nor NOR2_474 (G1729gat, G1694gat, G1695gat);
nor NOR2_475 (G1732gat, G1696gat, G1697gat);
nor NOR2_476 (G1735gat, G1698gat, G1699gat);
nor NOR2_477 (G1738gat, G1700gat, G1701gat);
nor NOR2_478 (G1741gat, G1702gat, G1703gat);
nor NOR2_479 (G1744gat, G1704gat, G1705gat);
nor NOR2_480 (G1747gat, G1706gat, G1707gat);
nor NOR2_481 (G1750gat, G1708gat, G1709gat);
nor NOR2_482 (G1753gat, G1710gat, G1711gat);
nor NOR2_483 (G1756gat, G1712gat, G1713gat);
nor NOR2_484 (G1759gat, G1714gat, G1221gat);
nor NOR2_485 (G1763gat, G1717gat, G549gat);
nor NOR2_486 (G1767gat, G1720gat, G597gat);
nor NOR2_487 (G1771gat, G1723gat, G645gat);
nor NOR2_488 (G1775gat, G1726gat, G693gat);
nor NOR2_489 (G1779gat, G1729gat, G741gat);
nor NOR2_490 (G1783gat, G1732gat, G789gat);
nor NOR2_491 (G1787gat, G1735gat, G837gat);
nor NOR2_492 (G1791gat, G1738gat, G885gat);
nor NOR2_493 (G1795gat, G1741gat, G933gat);
nor NOR2_494 (G1799gat, G1744gat, G981gat);
nor NOR2_495 (G1803gat, G1747gat, G1029gat);
nor NOR2_496 (G1807gat, G1750gat, G1077gat);
nor NOR2_497 (G1811gat, G1753gat, G1125gat);
nor NOR2_498 (G1815gat, G1756gat, G1173gat);
nor NOR2_499 (G1819gat, G1714gat, G1759gat);
nor NOR2_500 (G1820gat, G1759gat, G1221gat);
nor NOR2_501 (G1821gat, G1624gat, G1759gat);
nor NOR2_502 (G1824gat, G1717gat, G1763gat);
nor NOR2_503 (G1825gat, G1763gat, G549gat);
nor NOR2_504 (G1826gat, G1628gat, G1763gat);
nor NOR2_505 (G1829gat, G1720gat, G1767gat);
nor NOR2_506 (G1830gat, G1767gat, G597gat);
nor NOR2_507 (G1831gat, G1632gat, G1767gat);
nor NOR2_508 (G1834gat, G1723gat, G1771gat);
nor NOR2_509 (G1835gat, G1771gat, G645gat);
nor NOR2_510 (G1836gat, G1636gat, G1771gat);
nor NOR2_511 (G1839gat, G1726gat, G1775gat);
nor NOR2_512 (G1840gat, G1775gat, G693gat);
nor NOR2_513 (G1841gat, G1640gat, G1775gat);
nor NOR2_514 (G1844gat, G1729gat, G1779gat);
nor NOR2_515 (G1845gat, G1779gat, G741gat);
nor NOR2_516 (G1846gat, G1644gat, G1779gat);
nor NOR2_517 (G1849gat, G1732gat, G1783gat);
nor NOR2_518 (G1850gat, G1783gat, G789gat);
nor NOR2_519 (G1851gat, G1648gat, G1783gat);
nor NOR2_520 (G1854gat, G1735gat, G1787gat);
nor NOR2_521 (G1855gat, G1787gat, G837gat);
nor NOR2_522 (G1856gat, G1652gat, G1787gat);
nor NOR2_523 (G1859gat, G1738gat, G1791gat);
nor NOR2_524 (G1860gat, G1791gat, G885gat);
nor NOR2_525 (G1861gat, G1656gat, G1791gat);
nor NOR2_526 (G1864gat, G1741gat, G1795gat);
nor NOR2_527 (G1865gat, G1795gat, G933gat);
nor NOR2_528 (G1866gat, G1660gat, G1795gat);
nor NOR2_529 (G1869gat, G1744gat, G1799gat);
nor NOR2_530 (G1870gat, G1799gat, G981gat);
nor NOR2_531 (G1871gat, G1664gat, G1799gat);
nor NOR2_532 (G1874gat, G1747gat, G1803gat);
nor NOR2_533 (G1875gat, G1803gat, G1029gat);
nor NOR2_534 (G1876gat, G1668gat, G1803gat);
nor NOR2_535 (G1879gat, G1750gat, G1807gat);
nor NOR2_536 (G1880gat, G1807gat, G1077gat);
nor NOR2_537 (G1881gat, G1672gat, G1807gat);
nor NOR2_538 (G1884gat, G1753gat, G1811gat);
nor NOR2_539 (G1885gat, G1811gat, G1125gat);
nor NOR2_540 (G1886gat, G1676gat, G1811gat);
nor NOR2_541 (G1889gat, G1756gat, G1815gat);
nor NOR2_542 (G1890gat, G1815gat, G1173gat);
nor NOR2_543 (G1891gat, G1680gat, G1815gat);
nor NOR2_544 (G1894gat, G1819gat, G1820gat);
nor NOR2_545 (G1897gat, G1269gat, G1821gat);
nor NOR2_546 (G1901gat, G1824gat, G1825gat);
nor NOR2_547 (G1902gat, G1829gat, G1830gat);
nor NOR2_548 (G1905gat, G1834gat, G1835gat);
nor NOR2_549 (G1908gat, G1839gat, G1840gat);
nor NOR2_550 (G1911gat, G1844gat, G1845gat);
nor NOR2_551 (G1914gat, G1849gat, G1850gat);
nor NOR2_552 (G1917gat, G1854gat, G1855gat);
nor NOR2_553 (G1920gat, G1859gat, G1860gat);
nor NOR2_554 (G1923gat, G1864gat, G1865gat);
nor NOR2_555 (G1926gat, G1869gat, G1870gat);
nor NOR2_556 (G1929gat, G1874gat, G1875gat);
nor NOR2_557 (G1932gat, G1879gat, G1880gat);
nor NOR2_558 (G1935gat, G1884gat, G1885gat);
nor NOR2_559 (G1938gat, G1889gat, G1890gat);
nor NOR2_560 (G1941gat, G1894gat, G1891gat);
nor NOR2_561 (G1945gat, G1269gat, G1897gat);
nor NOR2_562 (G1946gat, G1897gat, G1821gat);
nor NOR2_563 (G1947gat, G1902gat, G1826gat);
nor NOR2_564 (G1951gat, G1905gat, G1831gat);
nor NOR2_565 (G1955gat, G1908gat, G1836gat);
nor NOR2_566 (G1959gat, G1911gat, G1841gat);
nor NOR2_567 (G1963gat, G1914gat, G1846gat);
nor NOR2_568 (G1967gat, G1917gat, G1851gat);
nor NOR2_569 (G1971gat, G1920gat, G1856gat);
nor NOR2_570 (G1975gat, G1923gat, G1861gat);
nor NOR2_571 (G1979gat, G1926gat, G1866gat);
nor NOR2_572 (G1983gat, G1929gat, G1871gat);
nor NOR2_573 (G1987gat, G1932gat, G1876gat);
nor NOR2_574 (G1991gat, G1935gat, G1881gat);
nor NOR2_575 (G1995gat, G1938gat, G1886gat);
nor NOR2_576 (G1999gat, G1894gat, G1941gat);
nor NOR2_577 (G2000gat, G1941gat, G1891gat);
nor NOR2_578 (G2001gat, G1945gat, G1946gat);
nor NOR2_579 (G2004gat, G1902gat, G1947gat);
nor NOR2_580 (G2005gat, G1947gat, G1826gat);
nor NOR2_581 (G2006gat, G1905gat, G1951gat);
nor NOR2_582 (G2007gat, G1951gat, G1831gat);
nor NOR2_583 (G2008gat, G1908gat, G1955gat);
nor NOR2_584 (G2009gat, G1955gat, G1836gat);
nor NOR2_585 (G2010gat, G1911gat, G1959gat);
nor NOR2_586 (G2011gat, G1959gat, G1841gat);
nor NOR2_587 (G2012gat, G1914gat, G1963gat);
nor NOR2_588 (G2013gat, G1963gat, G1846gat);
nor NOR2_589 (G2014gat, G1917gat, G1967gat);
nor NOR2_590 (G2015gat, G1967gat, G1851gat);
nor NOR2_591 (G2016gat, G1920gat, G1971gat);
nor NOR2_592 (G2017gat, G1971gat, G1856gat);
nor NOR2_593 (G2018gat, G1923gat, G1975gat);
nor NOR2_594 (G2019gat, G1975gat, G1861gat);
nor NOR2_595 (G2020gat, G1926gat, G1979gat);
nor NOR2_596 (G2021gat, G1979gat, G1866gat);
nor NOR2_597 (G2022gat, G1929gat, G1983gat);
nor NOR2_598 (G2023gat, G1983gat, G1871gat);
nor NOR2_599 (G2024gat, G1932gat, G1987gat);
nor NOR2_600 (G2025gat, G1987gat, G1876gat);
nor NOR2_601 (G2026gat, G1935gat, G1991gat);
nor NOR2_602 (G2027gat, G1991gat, G1881gat);
nor NOR2_603 (G2028gat, G1938gat, G1995gat);
nor NOR2_604 (G2029gat, G1995gat, G1886gat);
nor NOR2_605 (G2030gat, G1999gat, G2000gat);
nor NOR2_606 (G2033gat, G2001gat, G1224gat);
nor NOR2_607 (G2037gat, G2004gat, G2005gat);
nor NOR2_608 (G2040gat, G2006gat, G2007gat);
nor NOR2_609 (G2043gat, G2008gat, G2009gat);
nor NOR2_610 (G2046gat, G2010gat, G2011gat);
nor NOR2_611 (G2049gat, G2012gat, G2013gat);
nor NOR2_612 (G2052gat, G2014gat, G2015gat);
nor NOR2_613 (G2055gat, G2016gat, G2017gat);
nor NOR2_614 (G2058gat, G2018gat, G2019gat);
nor NOR2_615 (G2061gat, G2020gat, G2021gat);
nor NOR2_616 (G2064gat, G2022gat, G2023gat);
nor NOR2_617 (G2067gat, G2024gat, G2025gat);
nor NOR2_618 (G2070gat, G2026gat, G2027gat);
nor NOR2_619 (G2073gat, G2028gat, G2029gat);
nor NOR2_620 (G2076gat, G2030gat, G1176gat);
nor NOR2_621 (G2080gat, G2001gat, G2033gat);
nor NOR2_622 (G2081gat, G2033gat, G1224gat);
nor NOR2_623 (G2082gat, G1897gat, G2033gat);
nor NOR2_624 (G2085gat, G2037gat, G552gat);
nor NOR2_625 (G2089gat, G2040gat, G600gat);
nor NOR2_626 (G2093gat, G2043gat, G648gat);
nor NOR2_627 (G2097gat, G2046gat, G696gat);
nor NOR2_628 (G2101gat, G2049gat, G744gat);
nor NOR2_629 (G2105gat, G2052gat, G792gat);
nor NOR2_630 (G2109gat, G2055gat, G840gat);
nor NOR2_631 (G2113gat, G2058gat, G888gat);
nor NOR2_632 (G2117gat, G2061gat, G936gat);
nor NOR2_633 (G2121gat, G2064gat, G984gat);
nor NOR2_634 (G2125gat, G2067gat, G1032gat);
nor NOR2_635 (G2129gat, G2070gat, G1080gat);
nor NOR2_636 (G2133gat, G2073gat, G1128gat);
nor NOR2_637 (G2137gat, G2030gat, G2076gat);
nor NOR2_638 (G2138gat, G2076gat, G1176gat);
nor NOR2_639 (G2139gat, G1941gat, G2076gat);
nor NOR2_640 (G2142gat, G2080gat, G2081gat);
nor NOR2_641 (G2145gat, G1272gat, G2082gat);
nor NOR2_642 (G2149gat, G2037gat, G2085gat);
nor NOR2_643 (G2150gat, G2085gat, G552gat);
nor NOR2_644 (G2151gat, G1947gat, G2085gat);
nor NOR2_645 (G2154gat, G2040gat, G2089gat);
nor NOR2_646 (G2155gat, G2089gat, G600gat);
nor NOR2_647 (G2156gat, G1951gat, G2089gat);
nor NOR2_648 (G2159gat, G2043gat, G2093gat);
nor NOR2_649 (G2160gat, G2093gat, G648gat);
nor NOR2_650 (G2161gat, G1955gat, G2093gat);
nor NOR2_651 (G2164gat, G2046gat, G2097gat);
nor NOR2_652 (G2165gat, G2097gat, G696gat);
nor NOR2_653 (G2166gat, G1959gat, G2097gat);
nor NOR2_654 (G2169gat, G2049gat, G2101gat);
nor NOR2_655 (G2170gat, G2101gat, G744gat);
nor NOR2_656 (G2171gat, G1963gat, G2101gat);
nor NOR2_657 (G2174gat, G2052gat, G2105gat);
nor NOR2_658 (G2175gat, G2105gat, G792gat);
nor NOR2_659 (G2176gat, G1967gat, G2105gat);
nor NOR2_660 (G2179gat, G2055gat, G2109gat);
nor NOR2_661 (G2180gat, G2109gat, G840gat);
nor NOR2_662 (G2181gat, G1971gat, G2109gat);
nor NOR2_663 (G2184gat, G2058gat, G2113gat);
nor NOR2_664 (G2185gat, G2113gat, G888gat);
nor NOR2_665 (G2186gat, G1975gat, G2113gat);
nor NOR2_666 (G2189gat, G2061gat, G2117gat);
nor NOR2_667 (G2190gat, G2117gat, G936gat);
nor NOR2_668 (G2191gat, G1979gat, G2117gat);
nor NOR2_669 (G2194gat, G2064gat, G2121gat);
nor NOR2_670 (G2195gat, G2121gat, G984gat);
nor NOR2_671 (G2196gat, G1983gat, G2121gat);
nor NOR2_672 (G2199gat, G2067gat, G2125gat);
nor NOR2_673 (G2200gat, G2125gat, G1032gat);
nor NOR2_674 (G2201gat, G1987gat, G2125gat);
nor NOR2_675 (G2204gat, G2070gat, G2129gat);
nor NOR2_676 (G2205gat, G2129gat, G1080gat);
nor NOR2_677 (G2206gat, G1991gat, G2129gat);
nor NOR2_678 (G2209gat, G2073gat, G2133gat);
nor NOR2_679 (G2210gat, G2133gat, G1128gat);
nor NOR2_680 (G2211gat, G1995gat, G2133gat);
nor NOR2_681 (G2214gat, G2137gat, G2138gat);
nor NOR2_682 (G2217gat, G2142gat, G2139gat);
nor NOR2_683 (G2221gat, G1272gat, G2145gat);
nor NOR2_684 (G2222gat, G2145gat, G2082gat);
nor NOR2_685 (G2223gat, G2149gat, G2150gat);
nor NOR2_686 (G2224gat, G2154gat, G2155gat);
nor NOR2_687 (G2227gat, G2159gat, G2160gat);
nor NOR2_688 (G2230gat, G2164gat, G2165gat);
nor NOR2_689 (G2233gat, G2169gat, G2170gat);
nor NOR2_690 (G2236gat, G2174gat, G2175gat);
nor NOR2_691 (G2239gat, G2179gat, G2180gat);
nor NOR2_692 (G2242gat, G2184gat, G2185gat);
nor NOR2_693 (G2245gat, G2189gat, G2190gat);
nor NOR2_694 (G2248gat, G2194gat, G2195gat);
nor NOR2_695 (G2251gat, G2199gat, G2200gat);
nor NOR2_696 (G2254gat, G2204gat, G2205gat);
nor NOR2_697 (G2257gat, G2209gat, G2210gat);
nor NOR2_698 (G2260gat, G2214gat, G2211gat);
nor NOR2_699 (G2264gat, G2142gat, G2217gat);
nor NOR2_700 (G2265gat, G2217gat, G2139gat);
nor NOR2_701 (G2266gat, G2221gat, G2222gat);
nor NOR2_702 (G2269gat, G2224gat, G2151gat);
nor NOR2_703 (G2273gat, G2227gat, G2156gat);
nor NOR2_704 (G2277gat, G2230gat, G2161gat);
nor NOR2_705 (G2281gat, G2233gat, G2166gat);
nor NOR2_706 (G2285gat, G2236gat, G2171gat);
nor NOR2_707 (G2289gat, G2239gat, G2176gat);
nor NOR2_708 (G2293gat, G2242gat, G2181gat);
nor NOR2_709 (G2297gat, G2245gat, G2186gat);
nor NOR2_710 (G2301gat, G2248gat, G2191gat);
nor NOR2_711 (G2305gat, G2251gat, G2196gat);
nor NOR2_712 (G2309gat, G2254gat, G2201gat);
nor NOR2_713 (G2313gat, G2257gat, G2206gat);
nor NOR2_714 (G2317gat, G2214gat, G2260gat);
nor NOR2_715 (G2318gat, G2260gat, G2211gat);
nor NOR2_716 (G2319gat, G2264gat, G2265gat);
nor NOR2_717 (G2322gat, G2266gat, G1227gat);
nor NOR2_718 (G2326gat, G2224gat, G2269gat);
nor NOR2_719 (G2327gat, G2269gat, G2151gat);
nor NOR2_720 (G2328gat, G2227gat, G2273gat);
nor NOR2_721 (G2329gat, G2273gat, G2156gat);
nor NOR2_722 (G2330gat, G2230gat, G2277gat);
nor NOR2_723 (G2331gat, G2277gat, G2161gat);
nor NOR2_724 (G2332gat, G2233gat, G2281gat);
nor NOR2_725 (G2333gat, G2281gat, G2166gat);
nor NOR2_726 (G2334gat, G2236gat, G2285gat);
nor NOR2_727 (G2335gat, G2285gat, G2171gat);
nor NOR2_728 (G2336gat, G2239gat, G2289gat);
nor NOR2_729 (G2337gat, G2289gat, G2176gat);
nor NOR2_730 (G2338gat, G2242gat, G2293gat);
nor NOR2_731 (G2339gat, G2293gat, G2181gat);
nor NOR2_732 (G2340gat, G2245gat, G2297gat);
nor NOR2_733 (G2341gat, G2297gat, G2186gat);
nor NOR2_734 (G2342gat, G2248gat, G2301gat);
nor NOR2_735 (G2343gat, G2301gat, G2191gat);
nor NOR2_736 (G2344gat, G2251gat, G2305gat);
nor NOR2_737 (G2345gat, G2305gat, G2196gat);
nor NOR2_738 (G2346gat, G2254gat, G2309gat);
nor NOR2_739 (G2347gat, G2309gat, G2201gat);
nor NOR2_740 (G2348gat, G2257gat, G2313gat);
nor NOR2_741 (G2349gat, G2313gat, G2206gat);
nor NOR2_742 (G2350gat, G2317gat, G2318gat);
nor NOR2_743 (G2353gat, G2319gat, G1179gat);
nor NOR2_744 (G2357gat, G2266gat, G2322gat);
nor NOR2_745 (G2358gat, G2322gat, G1227gat);
nor NOR2_746 (G2359gat, G2145gat, G2322gat);
nor NOR2_747 (G2362gat, G2326gat, G2327gat);
nor NOR2_748 (G2365gat, G2328gat, G2329gat);
nor NOR2_749 (G2368gat, G2330gat, G2331gat);
nor NOR2_750 (G2371gat, G2332gat, G2333gat);
nor NOR2_751 (G2374gat, G2334gat, G2335gat);
nor NOR2_752 (G2377gat, G2336gat, G2337gat);
nor NOR2_753 (G2380gat, G2338gat, G2339gat);
nor NOR2_754 (G2383gat, G2340gat, G2341gat);
nor NOR2_755 (G2386gat, G2342gat, G2343gat);
nor NOR2_756 (G2389gat, G2344gat, G2345gat);
nor NOR2_757 (G2392gat, G2346gat, G2347gat);
nor NOR2_758 (G2395gat, G2348gat, G2349gat);
nor NOR2_759 (G2398gat, G2350gat, G1131gat);
nor NOR2_760 (G2402gat, G2319gat, G2353gat);
nor NOR2_761 (G2403gat, G2353gat, G1179gat);
nor NOR2_762 (G2404gat, G2217gat, G2353gat);
nor NOR2_763 (G2407gat, G2357gat, G2358gat);
nor NOR2_764 (G2410gat, G1275gat, G2359gat);
nor NOR2_765 (G2414gat, G2362gat, G555gat);
nor NOR2_766 (G2418gat, G2365gat, G603gat);
nor NOR2_767 (G2422gat, G2368gat, G651gat);
nor NOR2_768 (G2426gat, G2371gat, G699gat);
nor NOR2_769 (G2430gat, G2374gat, G747gat);
nor NOR2_770 (G2434gat, G2377gat, G795gat);
nor NOR2_771 (G2438gat, G2380gat, G843gat);
nor NOR2_772 (G2442gat, G2383gat, G891gat);
nor NOR2_773 (G2446gat, G2386gat, G939gat);
nor NOR2_774 (G2450gat, G2389gat, G987gat);
nor NOR2_775 (G2454gat, G2392gat, G1035gat);
nor NOR2_776 (G2458gat, G2395gat, G1083gat);
nor NOR2_777 (G2462gat, G2350gat, G2398gat);
nor NOR2_778 (G2463gat, G2398gat, G1131gat);
nor NOR2_779 (G2464gat, G2260gat, G2398gat);
nor NOR2_780 (G2467gat, G2402gat, G2403gat);
nor NOR2_781 (G2470gat, G2407gat, G2404gat);
nor NOR2_782 (G2474gat, G1275gat, G2410gat);
nor NOR2_783 (G2475gat, G2410gat, G2359gat);
nor NOR2_784 (G2476gat, G2362gat, G2414gat);
nor NOR2_785 (G2477gat, G2414gat, G555gat);
nor NOR2_786 (G2478gat, G2269gat, G2414gat);
nor NOR2_787 (G2481gat, G2365gat, G2418gat);
nor NOR2_788 (G2482gat, G2418gat, G603gat);
nor NOR2_789 (G2483gat, G2273gat, G2418gat);
nor NOR2_790 (G2486gat, G2368gat, G2422gat);
nor NOR2_791 (G2487gat, G2422gat, G651gat);
nor NOR2_792 (G2488gat, G2277gat, G2422gat);
nor NOR2_793 (G2491gat, G2371gat, G2426gat);
nor NOR2_794 (G2492gat, G2426gat, G699gat);
nor NOR2_795 (G2493gat, G2281gat, G2426gat);
nor NOR2_796 (G2496gat, G2374gat, G2430gat);
nor NOR2_797 (G2497gat, G2430gat, G747gat);
nor NOR2_798 (G2498gat, G2285gat, G2430gat);
nor NOR2_799 (G2501gat, G2377gat, G2434gat);
nor NOR2_800 (G2502gat, G2434gat, G795gat);
nor NOR2_801 (G2503gat, G2289gat, G2434gat);
nor NOR2_802 (G2506gat, G2380gat, G2438gat);
nor NOR2_803 (G2507gat, G2438gat, G843gat);
nor NOR2_804 (G2508gat, G2293gat, G2438gat);
nor NOR2_805 (G2511gat, G2383gat, G2442gat);
nor NOR2_806 (G2512gat, G2442gat, G891gat);
nor NOR2_807 (G2513gat, G2297gat, G2442gat);
nor NOR2_808 (G2516gat, G2386gat, G2446gat);
nor NOR2_809 (G2517gat, G2446gat, G939gat);
nor NOR2_810 (G2518gat, G2301gat, G2446gat);
nor NOR2_811 (G2521gat, G2389gat, G2450gat);
nor NOR2_812 (G2522gat, G2450gat, G987gat);
nor NOR2_813 (G2523gat, G2305gat, G2450gat);
nor NOR2_814 (G2526gat, G2392gat, G2454gat);
nor NOR2_815 (G2527gat, G2454gat, G1035gat);
nor NOR2_816 (G2528gat, G2309gat, G2454gat);
nor NOR2_817 (G2531gat, G2395gat, G2458gat);
nor NOR2_818 (G2532gat, G2458gat, G1083gat);
nor NOR2_819 (G2533gat, G2313gat, G2458gat);
nor NOR2_820 (G2536gat, G2462gat, G2463gat);
nor NOR2_821 (G2539gat, G2467gat, G2464gat);
nor NOR2_822 (G2543gat, G2407gat, G2470gat);
nor NOR2_823 (G2544gat, G2470gat, G2404gat);
nor NOR2_824 (G2545gat, G2474gat, G2475gat);
nor NOR2_825 (G2548gat, G2476gat, G2477gat);
nor NOR2_826 (G2549gat, G2481gat, G2482gat);
nor NOR2_827 (G2552gat, G2486gat, G2487gat);
nor NOR2_828 (G2555gat, G2491gat, G2492gat);
nor NOR2_829 (G2558gat, G2496gat, G2497gat);
nor NOR2_830 (G2561gat, G2501gat, G2502gat);
nor NOR2_831 (G2564gat, G2506gat, G2507gat);
nor NOR2_832 (G2567gat, G2511gat, G2512gat);
nor NOR2_833 (G2570gat, G2516gat, G2517gat);
nor NOR2_834 (G2573gat, G2521gat, G2522gat);
nor NOR2_835 (G2576gat, G2526gat, G2527gat);
nor NOR2_836 (G2579gat, G2531gat, G2532gat);
nor NOR2_837 (G2582gat, G2536gat, G2533gat);
nor NOR2_838 (G2586gat, G2467gat, G2539gat);
nor NOR2_839 (G2587gat, G2539gat, G2464gat);
nor NOR2_840 (G2588gat, G2543gat, G2544gat);
nor NOR2_841 (G2591gat, G2545gat, G1230gat);
nor NOR2_842 (G2595gat, G2549gat, G2478gat);
nor NOR2_843 (G2599gat, G2552gat, G2483gat);
nor NOR2_844 (G2603gat, G2555gat, G2488gat);
nor NOR2_845 (G2607gat, G2558gat, G2493gat);
nor NOR2_846 (G2611gat, G2561gat, G2498gat);
nor NOR2_847 (G2615gat, G2564gat, G2503gat);
nor NOR2_848 (G2619gat, G2567gat, G2508gat);
nor NOR2_849 (G2623gat, G2570gat, G2513gat);
nor NOR2_850 (G2627gat, G2573gat, G2518gat);
nor NOR2_851 (G2631gat, G2576gat, G2523gat);
nor NOR2_852 (G2635gat, G2579gat, G2528gat);
nor NOR2_853 (G2639gat, G2536gat, G2582gat);
nor NOR2_854 (G2640gat, G2582gat, G2533gat);
nor NOR2_855 (G2641gat, G2586gat, G2587gat);
nor NOR2_856 (G2644gat, G2588gat, G1182gat);
nor NOR2_857 (G2648gat, G2545gat, G2591gat);
nor NOR2_858 (G2649gat, G2591gat, G1230gat);
nor NOR2_859 (G2650gat, G2410gat, G2591gat);
nor NOR2_860 (G2653gat, G2549gat, G2595gat);
nor NOR2_861 (G2654gat, G2595gat, G2478gat);
nor NOR2_862 (G2655gat, G2552gat, G2599gat);
nor NOR2_863 (G2656gat, G2599gat, G2483gat);
nor NOR2_864 (G2657gat, G2555gat, G2603gat);
nor NOR2_865 (G2658gat, G2603gat, G2488gat);
nor NOR2_866 (G2659gat, G2558gat, G2607gat);
nor NOR2_867 (G2660gat, G2607gat, G2493gat);
nor NOR2_868 (G2661gat, G2561gat, G2611gat);
nor NOR2_869 (G2662gat, G2611gat, G2498gat);
nor NOR2_870 (G2663gat, G2564gat, G2615gat);
nor NOR2_871 (G2664gat, G2615gat, G2503gat);
nor NOR2_872 (G2665gat, G2567gat, G2619gat);
nor NOR2_873 (G2666gat, G2619gat, G2508gat);
nor NOR2_874 (G2667gat, G2570gat, G2623gat);
nor NOR2_875 (G2668gat, G2623gat, G2513gat);
nor NOR2_876 (G2669gat, G2573gat, G2627gat);
nor NOR2_877 (G2670gat, G2627gat, G2518gat);
nor NOR2_878 (G2671gat, G2576gat, G2631gat);
nor NOR2_879 (G2672gat, G2631gat, G2523gat);
nor NOR2_880 (G2673gat, G2579gat, G2635gat);
nor NOR2_881 (G2674gat, G2635gat, G2528gat);
nor NOR2_882 (G2675gat, G2639gat, G2640gat);
nor NOR2_883 (G2678gat, G2641gat, G1134gat);
nor NOR2_884 (G2682gat, G2588gat, G2644gat);
nor NOR2_885 (G2683gat, G2644gat, G1182gat);
nor NOR2_886 (G2684gat, G2470gat, G2644gat);
nor NOR2_887 (G2687gat, G2648gat, G2649gat);
nor NOR2_888 (G2690gat, G1278gat, G2650gat);
nor NOR2_889 (G2694gat, G2653gat, G2654gat);
nor NOR2_890 (G2697gat, G2655gat, G2656gat);
nor NOR2_891 (G2700gat, G2657gat, G2658gat);
nor NOR2_892 (G2703gat, G2659gat, G2660gat);
nor NOR2_893 (G2706gat, G2661gat, G2662gat);
nor NOR2_894 (G2709gat, G2663gat, G2664gat);
nor NOR2_895 (G2712gat, G2665gat, G2666gat);
nor NOR2_896 (G2715gat, G2667gat, G2668gat);
nor NOR2_897 (G2718gat, G2669gat, G2670gat);
nor NOR2_898 (G2721gat, G2671gat, G2672gat);
nor NOR2_899 (G2724gat, G2673gat, G2674gat);
nor NOR2_900 (G2727gat, G2675gat, G1086gat);
nor NOR2_901 (G2731gat, G2641gat, G2678gat);
nor NOR2_902 (G2732gat, G2678gat, G1134gat);
nor NOR2_903 (G2733gat, G2539gat, G2678gat);
nor NOR2_904 (G2736gat, G2682gat, G2683gat);
nor NOR2_905 (G2739gat, G2687gat, G2684gat);
nor NOR2_906 (G2743gat, G1278gat, G2690gat);
nor NOR2_907 (G2744gat, G2690gat, G2650gat);
nor NOR2_908 (G2745gat, G2694gat, G558gat);
nor NOR2_909 (G2749gat, G2697gat, G606gat);
nor NOR2_910 (G2753gat, G2700gat, G654gat);
nor NOR2_911 (G2757gat, G2703gat, G702gat);
nor NOR2_912 (G2761gat, G2706gat, G750gat);
nor NOR2_913 (G2765gat, G2709gat, G798gat);
nor NOR2_914 (G2769gat, G2712gat, G846gat);
nor NOR2_915 (G2773gat, G2715gat, G894gat);
nor NOR2_916 (G2777gat, G2718gat, G942gat);
nor NOR2_917 (G2781gat, G2721gat, G990gat);
nor NOR2_918 (G2785gat, G2724gat, G1038gat);
nor NOR2_919 (G2789gat, G2675gat, G2727gat);
nor NOR2_920 (G2790gat, G2727gat, G1086gat);
nor NOR2_921 (G2791gat, G2582gat, G2727gat);
nor NOR2_922 (G2794gat, G2731gat, G2732gat);
nor NOR2_923 (G2797gat, G2736gat, G2733gat);
nor NOR2_924 (G2801gat, G2687gat, G2739gat);
nor NOR2_925 (G2802gat, G2739gat, G2684gat);
nor NOR2_926 (G2803gat, G2743gat, G2744gat);
nor NOR2_927 (G2806gat, G2694gat, G2745gat);
nor NOR2_928 (G2807gat, G2745gat, G558gat);
nor NOR2_929 (G2808gat, G2595gat, G2745gat);
nor NOR2_930 (G2811gat, G2697gat, G2749gat);
nor NOR2_931 (G2812gat, G2749gat, G606gat);
nor NOR2_932 (G2813gat, G2599gat, G2749gat);
nor NOR2_933 (G2816gat, G2700gat, G2753gat);
nor NOR2_934 (G2817gat, G2753gat, G654gat);
nor NOR2_935 (G2818gat, G2603gat, G2753gat);
nor NOR2_936 (G2821gat, G2703gat, G2757gat);
nor NOR2_937 (G2822gat, G2757gat, G702gat);
nor NOR2_938 (G2823gat, G2607gat, G2757gat);
nor NOR2_939 (G2826gat, G2706gat, G2761gat);
nor NOR2_940 (G2827gat, G2761gat, G750gat);
nor NOR2_941 (G2828gat, G2611gat, G2761gat);
nor NOR2_942 (G2831gat, G2709gat, G2765gat);
nor NOR2_943 (G2832gat, G2765gat, G798gat);
nor NOR2_944 (G2833gat, G2615gat, G2765gat);
nor NOR2_945 (G2836gat, G2712gat, G2769gat);
nor NOR2_946 (G2837gat, G2769gat, G846gat);
nor NOR2_947 (G2838gat, G2619gat, G2769gat);
nor NOR2_948 (G2841gat, G2715gat, G2773gat);
nor NOR2_949 (G2842gat, G2773gat, G894gat);
nor NOR2_950 (G2843gat, G2623gat, G2773gat);
nor NOR2_951 (G2846gat, G2718gat, G2777gat);
nor NOR2_952 (G2847gat, G2777gat, G942gat);
nor NOR2_953 (G2848gat, G2627gat, G2777gat);
nor NOR2_954 (G2851gat, G2721gat, G2781gat);
nor NOR2_955 (G2852gat, G2781gat, G990gat);
nor NOR2_956 (G2853gat, G2631gat, G2781gat);
nor NOR2_957 (G2856gat, G2724gat, G2785gat);
nor NOR2_958 (G2857gat, G2785gat, G1038gat);
nor NOR2_959 (G2858gat, G2635gat, G2785gat);
nor NOR2_960 (G2861gat, G2789gat, G2790gat);
nor NOR2_961 (G2864gat, G2794gat, G2791gat);
nor NOR2_962 (G2868gat, G2736gat, G2797gat);
nor NOR2_963 (G2869gat, G2797gat, G2733gat);
nor NOR2_964 (G2870gat, G2801gat, G2802gat);
nor NOR2_965 (G2873gat, G2803gat, G1233gat);
nor NOR2_966 (G2877gat, G2806gat, G2807gat);
nor NOR2_967 (G2878gat, G2811gat, G2812gat);
nor NOR2_968 (G2881gat, G2816gat, G2817gat);
nor NOR2_969 (G2884gat, G2821gat, G2822gat);
nor NOR2_970 (G2887gat, G2826gat, G2827gat);
nor NOR2_971 (G2890gat, G2831gat, G2832gat);
nor NOR2_972 (G2893gat, G2836gat, G2837gat);
nor NOR2_973 (G2896gat, G2841gat, G2842gat);
nor NOR2_974 (G2899gat, G2846gat, G2847gat);
nor NOR2_975 (G2902gat, G2851gat, G2852gat);
nor NOR2_976 (G2905gat, G2856gat, G2857gat);
nor NOR2_977 (G2908gat, G2861gat, G2858gat);
nor NOR2_978 (G2912gat, G2794gat, G2864gat);
nor NOR2_979 (G2913gat, G2864gat, G2791gat);
nor NOR2_980 (G2914gat, G2868gat, G2869gat);
nor NOR2_981 (G2917gat, G2870gat, G1185gat);
nor NOR2_982 (G2921gat, G2803gat, G2873gat);
nor NOR2_983 (G2922gat, G2873gat, G1233gat);
nor NOR2_984 (G2923gat, G2690gat, G2873gat);
nor NOR2_985 (G2926gat, G2878gat, G2808gat);
nor NOR2_986 (G2930gat, G2881gat, G2813gat);
nor NOR2_987 (G2934gat, G2884gat, G2818gat);
nor NOR2_988 (G2938gat, G2887gat, G2823gat);
nor NOR2_989 (G2942gat, G2890gat, G2828gat);
nor NOR2_990 (G2946gat, G2893gat, G2833gat);
nor NOR2_991 (G2950gat, G2896gat, G2838gat);
nor NOR2_992 (G2954gat, G2899gat, G2843gat);
nor NOR2_993 (G2958gat, G2902gat, G2848gat);
nor NOR2_994 (G2962gat, G2905gat, G2853gat);
nor NOR2_995 (G2966gat, G2861gat, G2908gat);
nor NOR2_996 (G2967gat, G2908gat, G2858gat);
nor NOR2_997 (G2968gat, G2912gat, G2913gat);
nor NOR2_998 (G2971gat, G2914gat, G1137gat);
nor NOR2_999 (G2975gat, G2870gat, G2917gat);
nor NOR2_1000 (G2976gat, G2917gat, G1185gat);
nor NOR2_1001 (G2977gat, G2739gat, G2917gat);
nor NOR2_1002 (G2980gat, G2921gat, G2922gat);
nor NOR2_1003 (G2983gat, G1281gat, G2923gat);
nor NOR2_1004 (G2987gat, G2878gat, G2926gat);
nor NOR2_1005 (G2988gat, G2926gat, G2808gat);
nor NOR2_1006 (G2989gat, G2881gat, G2930gat);
nor NOR2_1007 (G2990gat, G2930gat, G2813gat);
nor NOR2_1008 (G2991gat, G2884gat, G2934gat);
nor NOR2_1009 (G2992gat, G2934gat, G2818gat);
nor NOR2_1010 (G2993gat, G2887gat, G2938gat);
nor NOR2_1011 (G2994gat, G2938gat, G2823gat);
nor NOR2_1012 (G2995gat, G2890gat, G2942gat);
nor NOR2_1013 (G2996gat, G2942gat, G2828gat);
nor NOR2_1014 (G2997gat, G2893gat, G2946gat);
nor NOR2_1015 (G2998gat, G2946gat, G2833gat);
nor NOR2_1016 (G2999gat, G2896gat, G2950gat);
nor NOR2_1017 (G3000gat, G2950gat, G2838gat);
nor NOR2_1018 (G3001gat, G2899gat, G2954gat);
nor NOR2_1019 (G3002gat, G2954gat, G2843gat);
nor NOR2_1020 (G3003gat, G2902gat, G2958gat);
nor NOR2_1021 (G3004gat, G2958gat, G2848gat);
nor NOR2_1022 (G3005gat, G2905gat, G2962gat);
nor NOR2_1023 (G3006gat, G2962gat, G2853gat);
nor NOR2_1024 (G3007gat, G2966gat, G2967gat);
nor NOR2_1025 (G3010gat, G2968gat, G1089gat);
nor NOR2_1026 (G3014gat, G2914gat, G2971gat);
nor NOR2_1027 (G3015gat, G2971gat, G1137gat);
nor NOR2_1028 (G3016gat, G2797gat, G2971gat);
nor NOR2_1029 (G3019gat, G2975gat, G2976gat);
nor NOR2_1030 (G3022gat, G2980gat, G2977gat);
nor NOR2_1031 (G3026gat, G1281gat, G2983gat);
nor NOR2_1032 (G3027gat, G2983gat, G2923gat);
nor NOR2_1033 (G3028gat, G2987gat, G2988gat);
nor NOR2_1034 (G3031gat, G2989gat, G2990gat);
nor NOR2_1035 (G3034gat, G2991gat, G2992gat);
nor NOR2_1036 (G3037gat, G2993gat, G2994gat);
nor NOR2_1037 (G3040gat, G2995gat, G2996gat);
nor NOR2_1038 (G3043gat, G2997gat, G2998gat);
nor NOR2_1039 (G3046gat, G2999gat, G3000gat);
nor NOR2_1040 (G3049gat, G3001gat, G3002gat);
nor NOR2_1041 (G3052gat, G3003gat, G3004gat);
nor NOR2_1042 (G3055gat, G3005gat, G3006gat);
nor NOR2_1043 (G3058gat, G3007gat, G1041gat);
nor NOR2_1044 (G3062gat, G2968gat, G3010gat);
nor NOR2_1045 (G3063gat, G3010gat, G1089gat);
nor NOR2_1046 (G3064gat, G2864gat, G3010gat);
nor NOR2_1047 (G3067gat, G3014gat, G3015gat);
nor NOR2_1048 (G3070gat, G3019gat, G3016gat);
nor NOR2_1049 (G3074gat, G2980gat, G3022gat);
nor NOR2_1050 (G3075gat, G3022gat, G2977gat);
nor NOR2_1051 (G3076gat, G3026gat, G3027gat);
nor NOR2_1052 (G3079gat, G3028gat, G561gat);
nor NOR2_1053 (G3083gat, G3031gat, G609gat);
nor NOR2_1054 (G3087gat, G3034gat, G657gat);
nor NOR2_1055 (G3091gat, G3037gat, G705gat);
nor NOR2_1056 (G3095gat, G3040gat, G753gat);
nor NOR2_1057 (G3099gat, G3043gat, G801gat);
nor NOR2_1058 (G3103gat, G3046gat, G849gat);
nor NOR2_1059 (G3107gat, G3049gat, G897gat);
nor NOR2_1060 (G3111gat, G3052gat, G945gat);
nor NOR2_1061 (G3115gat, G3055gat, G993gat);
nor NOR2_1062 (G3119gat, G3007gat, G3058gat);
nor NOR2_1063 (G3120gat, G3058gat, G1041gat);
nor NOR2_1064 (G3121gat, G2908gat, G3058gat);
nor NOR2_1065 (G3124gat, G3062gat, G3063gat);
nor NOR2_1066 (G3127gat, G3067gat, G3064gat);
nor NOR2_1067 (G3131gat, G3019gat, G3070gat);
nor NOR2_1068 (G3132gat, G3070gat, G3016gat);
nor NOR2_1069 (G3133gat, G3074gat, G3075gat);
nor NOR2_1070 (G3136gat, G3076gat, G1236gat);
nor NOR2_1071 (G3140gat, G3028gat, G3079gat);
nor NOR2_1072 (G3141gat, G3079gat, G561gat);
nor NOR2_1073 (G3142gat, G2926gat, G3079gat);
nor NOR2_1074 (G3145gat, G3031gat, G3083gat);
nor NOR2_1075 (G3146gat, G3083gat, G609gat);
nor NOR2_1076 (G3147gat, G2930gat, G3083gat);
nor NOR2_1077 (G3150gat, G3034gat, G3087gat);
nor NOR2_1078 (G3151gat, G3087gat, G657gat);
nor NOR2_1079 (G3152gat, G2934gat, G3087gat);
nor NOR2_1080 (G3155gat, G3037gat, G3091gat);
nor NOR2_1081 (G3156gat, G3091gat, G705gat);
nor NOR2_1082 (G3157gat, G2938gat, G3091gat);
nor NOR2_1083 (G3160gat, G3040gat, G3095gat);
nor NOR2_1084 (G3161gat, G3095gat, G753gat);
nor NOR2_1085 (G3162gat, G2942gat, G3095gat);
nor NOR2_1086 (G3165gat, G3043gat, G3099gat);
nor NOR2_1087 (G3166gat, G3099gat, G801gat);
nor NOR2_1088 (G3167gat, G2946gat, G3099gat);
nor NOR2_1089 (G3170gat, G3046gat, G3103gat);
nor NOR2_1090 (G3171gat, G3103gat, G849gat);
nor NOR2_1091 (G3172gat, G2950gat, G3103gat);
nor NOR2_1092 (G3175gat, G3049gat, G3107gat);
nor NOR2_1093 (G3176gat, G3107gat, G897gat);
nor NOR2_1094 (G3177gat, G2954gat, G3107gat);
nor NOR2_1095 (G3180gat, G3052gat, G3111gat);
nor NOR2_1096 (G3181gat, G3111gat, G945gat);
nor NOR2_1097 (G3182gat, G2958gat, G3111gat);
nor NOR2_1098 (G3185gat, G3055gat, G3115gat);
nor NOR2_1099 (G3186gat, G3115gat, G993gat);
nor NOR2_1100 (G3187gat, G2962gat, G3115gat);
nor NOR2_1101 (G3190gat, G3119gat, G3120gat);
nor NOR2_1102 (G3193gat, G3124gat, G3121gat);
nor NOR2_1103 (G3197gat, G3067gat, G3127gat);
nor NOR2_1104 (G3198gat, G3127gat, G3064gat);
nor NOR2_1105 (G3199gat, G3131gat, G3132gat);
nor NOR2_1106 (G3202gat, G3133gat, G1188gat);
nor NOR2_1107 (G3206gat, G3076gat, G3136gat);
nor NOR2_1108 (G3207gat, G3136gat, G1236gat);
nor NOR2_1109 (G3208gat, G2983gat, G3136gat);
nor NOR2_1110 (G3211gat, G3140gat, G3141gat);
nor NOR2_1111 (G3212gat, G3145gat, G3146gat);
nor NOR2_1112 (G3215gat, G3150gat, G3151gat);
nor NOR2_1113 (G3218gat, G3155gat, G3156gat);
nor NOR2_1114 (G3221gat, G3160gat, G3161gat);
nor NOR2_1115 (G3224gat, G3165gat, G3166gat);
nor NOR2_1116 (G3227gat, G3170gat, G3171gat);
nor NOR2_1117 (G3230gat, G3175gat, G3176gat);
nor NOR2_1118 (G3233gat, G3180gat, G3181gat);
nor NOR2_1119 (G3236gat, G3185gat, G3186gat);
nor NOR2_1120 (G3239gat, G3190gat, G3187gat);
nor NOR2_1121 (G3243gat, G3124gat, G3193gat);
nor NOR2_1122 (G3244gat, G3193gat, G3121gat);
nor NOR2_1123 (G3245gat, G3197gat, G3198gat);
nor NOR2_1124 (G3248gat, G3199gat, G1140gat);
nor NOR2_1125 (G3252gat, G3133gat, G3202gat);
nor NOR2_1126 (G3253gat, G3202gat, G1188gat);
nor NOR2_1127 (G3254gat, G3022gat, G3202gat);
nor NOR2_1128 (G3257gat, G3206gat, G3207gat);
nor NOR2_1129 (G3260gat, G1284gat, G3208gat);
nor NOR2_1130 (G3264gat, G3212gat, G3142gat);
nor NOR2_1131 (G3268gat, G3215gat, G3147gat);
nor NOR2_1132 (G3272gat, G3218gat, G3152gat);
nor NOR2_1133 (G3276gat, G3221gat, G3157gat);
nor NOR2_1134 (G3280gat, G3224gat, G3162gat);
nor NOR2_1135 (G3284gat, G3227gat, G3167gat);
nor NOR2_1136 (G3288gat, G3230gat, G3172gat);
nor NOR2_1137 (G3292gat, G3233gat, G3177gat);
nor NOR2_1138 (G3296gat, G3236gat, G3182gat);
nor NOR2_1139 (G3300gat, G3190gat, G3239gat);
nor NOR2_1140 (G3301gat, G3239gat, G3187gat);
nor NOR2_1141 (G3302gat, G3243gat, G3244gat);
nor NOR2_1142 (G3305gat, G3245gat, G1092gat);
nor NOR2_1143 (G3309gat, G3199gat, G3248gat);
nor NOR2_1144 (G3310gat, G3248gat, G1140gat);
nor NOR2_1145 (G3311gat, G3070gat, G3248gat);
nor NOR2_1146 (G3314gat, G3252gat, G3253gat);
nor NOR2_1147 (G3317gat, G3257gat, G3254gat);
nor NOR2_1148 (G3321gat, G1284gat, G3260gat);
nor NOR2_1149 (G3322gat, G3260gat, G3208gat);
nor NOR2_1150 (G3323gat, G3212gat, G3264gat);
nor NOR2_1151 (G3324gat, G3264gat, G3142gat);
nor NOR2_1152 (G3325gat, G3215gat, G3268gat);
nor NOR2_1153 (G3326gat, G3268gat, G3147gat);
nor NOR2_1154 (G3327gat, G3218gat, G3272gat);
nor NOR2_1155 (G3328gat, G3272gat, G3152gat);
nor NOR2_1156 (G3329gat, G3221gat, G3276gat);
nor NOR2_1157 (G3330gat, G3276gat, G3157gat);
nor NOR2_1158 (G3331gat, G3224gat, G3280gat);
nor NOR2_1159 (G3332gat, G3280gat, G3162gat);
nor NOR2_1160 (G3333gat, G3227gat, G3284gat);
nor NOR2_1161 (G3334gat, G3284gat, G3167gat);
nor NOR2_1162 (G3335gat, G3230gat, G3288gat);
nor NOR2_1163 (G3336gat, G3288gat, G3172gat);
nor NOR2_1164 (G3337gat, G3233gat, G3292gat);
nor NOR2_1165 (G3338gat, G3292gat, G3177gat);
nor NOR2_1166 (G3339gat, G3236gat, G3296gat);
nor NOR2_1167 (G3340gat, G3296gat, G3182gat);
nor NOR2_1168 (G3341gat, G3300gat, G3301gat);
nor NOR2_1169 (G3344gat, G3302gat, G1044gat);
nor NOR2_1170 (G3348gat, G3245gat, G3305gat);
nor NOR2_1171 (G3349gat, G3305gat, G1092gat);
nor NOR2_1172 (G3350gat, G3127gat, G3305gat);
nor NOR2_1173 (G3353gat, G3309gat, G3310gat);
nor NOR2_1174 (G3356gat, G3314gat, G3311gat);
nor NOR2_1175 (G3360gat, G3257gat, G3317gat);
nor NOR2_1176 (G3361gat, G3317gat, G3254gat);
nor NOR2_1177 (G3362gat, G3321gat, G3322gat);
nor NOR2_1178 (G3365gat, G3323gat, G3324gat);
nor NOR2_1179 (G3368gat, G3325gat, G3326gat);
nor NOR2_1180 (G3371gat, G3327gat, G3328gat);
nor NOR2_1181 (G3374gat, G3329gat, G3330gat);
nor NOR2_1182 (G3377gat, G3331gat, G3332gat);
nor NOR2_1183 (G3380gat, G3333gat, G3334gat);
nor NOR2_1184 (G3383gat, G3335gat, G3336gat);
nor NOR2_1185 (G3386gat, G3337gat, G3338gat);
nor NOR2_1186 (G3389gat, G3339gat, G3340gat);
nor NOR2_1187 (G3392gat, G3341gat, G996gat);
nor NOR2_1188 (G3396gat, G3302gat, G3344gat);
nor NOR2_1189 (G3397gat, G3344gat, G1044gat);
nor NOR2_1190 (G3398gat, G3193gat, G3344gat);
nor NOR2_1191 (G3401gat, G3348gat, G3349gat);
nor NOR2_1192 (G3404gat, G3353gat, G3350gat);
nor NOR2_1193 (G3408gat, G3314gat, G3356gat);
nor NOR2_1194 (G3409gat, G3356gat, G3311gat);
nor NOR2_1195 (G3410gat, G3360gat, G3361gat);
nor NOR2_1196 (G3413gat, G3362gat, G1239gat);
nor NOR2_1197 (G3417gat, G3365gat, G564gat);
nor NOR2_1198 (G3421gat, G3368gat, G612gat);
nor NOR2_1199 (G3425gat, G3371gat, G660gat);
nor NOR2_1200 (G3429gat, G3374gat, G708gat);
nor NOR2_1201 (G3433gat, G3377gat, G756gat);
nor NOR2_1202 (G3437gat, G3380gat, G804gat);
nor NOR2_1203 (G3441gat, G3383gat, G852gat);
nor NOR2_1204 (G3445gat, G3386gat, G900gat);
nor NOR2_1205 (G3449gat, G3389gat, G948gat);
nor NOR2_1206 (G3453gat, G3341gat, G3392gat);
nor NOR2_1207 (G3454gat, G3392gat, G996gat);
nor NOR2_1208 (G3455gat, G3239gat, G3392gat);
nor NOR2_1209 (G3458gat, G3396gat, G3397gat);
nor NOR2_1210 (G3461gat, G3401gat, G3398gat);
nor NOR2_1211 (G3465gat, G3353gat, G3404gat);
nor NOR2_1212 (G3466gat, G3404gat, G3350gat);
nor NOR2_1213 (G3467gat, G3408gat, G3409gat);
nor NOR2_1214 (G3470gat, G3410gat, G1191gat);
nor NOR2_1215 (G3474gat, G3362gat, G3413gat);
nor NOR2_1216 (G3475gat, G3413gat, G1239gat);
nor NOR2_1217 (G3476gat, G3260gat, G3413gat);
nor NOR2_1218 (G3479gat, G3365gat, G3417gat);
nor NOR2_1219 (G3480gat, G3417gat, G564gat);
nor NOR2_1220 (G3481gat, G3264gat, G3417gat);
nor NOR2_1221 (G3484gat, G3368gat, G3421gat);
nor NOR2_1222 (G3485gat, G3421gat, G612gat);
nor NOR2_1223 (G3486gat, G3268gat, G3421gat);
nor NOR2_1224 (G3489gat, G3371gat, G3425gat);
nor NOR2_1225 (G3490gat, G3425gat, G660gat);
nor NOR2_1226 (G3491gat, G3272gat, G3425gat);
nor NOR2_1227 (G3494gat, G3374gat, G3429gat);
nor NOR2_1228 (G3495gat, G3429gat, G708gat);
nor NOR2_1229 (G3496gat, G3276gat, G3429gat);
nor NOR2_1230 (G3499gat, G3377gat, G3433gat);
nor NOR2_1231 (G3500gat, G3433gat, G756gat);
nor NOR2_1232 (G3501gat, G3280gat, G3433gat);
nor NOR2_1233 (G3504gat, G3380gat, G3437gat);
nor NOR2_1234 (G3505gat, G3437gat, G804gat);
nor NOR2_1235 (G3506gat, G3284gat, G3437gat);
nor NOR2_1236 (G3509gat, G3383gat, G3441gat);
nor NOR2_1237 (G3510gat, G3441gat, G852gat);
nor NOR2_1238 (G3511gat, G3288gat, G3441gat);
nor NOR2_1239 (G3514gat, G3386gat, G3445gat);
nor NOR2_1240 (G3515gat, G3445gat, G900gat);
nor NOR2_1241 (G3516gat, G3292gat, G3445gat);
nor NOR2_1242 (G3519gat, G3389gat, G3449gat);
nor NOR2_1243 (G3520gat, G3449gat, G948gat);
nor NOR2_1244 (G3521gat, G3296gat, G3449gat);
nor NOR2_1245 (G3524gat, G3453gat, G3454gat);
nor NOR2_1246 (G3527gat, G3458gat, G3455gat);
nor NOR2_1247 (G3531gat, G3401gat, G3461gat);
nor NOR2_1248 (G3532gat, G3461gat, G3398gat);
nor NOR2_1249 (G3533gat, G3465gat, G3466gat);
nor NOR2_1250 (G3536gat, G3467gat, G1143gat);
nor NOR2_1251 (G3540gat, G3410gat, G3470gat);
nor NOR2_1252 (G3541gat, G3470gat, G1191gat);
nor NOR2_1253 (G3542gat, G3317gat, G3470gat);
nor NOR2_1254 (G3545gat, G3474gat, G3475gat);
nor NOR2_1255 (G3548gat, G1287gat, G3476gat);
nor NOR2_1256 (G3552gat, G3479gat, G3480gat);
nor NOR2_1257 (G3553gat, G3484gat, G3485gat);
nor NOR2_1258 (G3556gat, G3489gat, G3490gat);
nor NOR2_1259 (G3559gat, G3494gat, G3495gat);
nor NOR2_1260 (G3562gat, G3499gat, G3500gat);
nor NOR2_1261 (G3565gat, G3504gat, G3505gat);
nor NOR2_1262 (G3568gat, G3509gat, G3510gat);
nor NOR2_1263 (G3571gat, G3514gat, G3515gat);
nor NOR2_1264 (G3574gat, G3519gat, G3520gat);
nor NOR2_1265 (G3577gat, G3524gat, G3521gat);
nor NOR2_1266 (G3581gat, G3458gat, G3527gat);
nor NOR2_1267 (G3582gat, G3527gat, G3455gat);
nor NOR2_1268 (G3583gat, G3531gat, G3532gat);
nor NOR2_1269 (G3586gat, G3533gat, G1095gat);
nor NOR2_1270 (G3590gat, G3467gat, G3536gat);
nor NOR2_1271 (G3591gat, G3536gat, G1143gat);
nor NOR2_1272 (G3592gat, G3356gat, G3536gat);
nor NOR2_1273 (G3595gat, G3540gat, G3541gat);
nor NOR2_1274 (G3598gat, G3545gat, G3542gat);
nor NOR2_1275 (G3602gat, G1287gat, G3548gat);
nor NOR2_1276 (G3603gat, G3548gat, G3476gat);
nor NOR2_1277 (G3604gat, G3553gat, G3481gat);
nor NOR2_1278 (G3608gat, G3556gat, G3486gat);
nor NOR2_1279 (G3612gat, G3559gat, G3491gat);
nor NOR2_1280 (G3616gat, G3562gat, G3496gat);
nor NOR2_1281 (G3620gat, G3565gat, G3501gat);
nor NOR2_1282 (G3624gat, G3568gat, G3506gat);
nor NOR2_1283 (G3628gat, G3571gat, G3511gat);
nor NOR2_1284 (G3632gat, G3574gat, G3516gat);
nor NOR2_1285 (G3636gat, G3524gat, G3577gat);
nor NOR2_1286 (G3637gat, G3577gat, G3521gat);
nor NOR2_1287 (G3638gat, G3581gat, G3582gat);
nor NOR2_1288 (G3641gat, G3583gat, G1047gat);
nor NOR2_1289 (G3645gat, G3533gat, G3586gat);
nor NOR2_1290 (G3646gat, G3586gat, G1095gat);
nor NOR2_1291 (G3647gat, G3404gat, G3586gat);
nor NOR2_1292 (G3650gat, G3590gat, G3591gat);
nor NOR2_1293 (G3653gat, G3595gat, G3592gat);
nor NOR2_1294 (G3657gat, G3545gat, G3598gat);
nor NOR2_1295 (G3658gat, G3598gat, G3542gat);
nor NOR2_1296 (G3659gat, G3602gat, G3603gat);
nor NOR2_1297 (G3662gat, G3553gat, G3604gat);
nor NOR2_1298 (G3663gat, G3604gat, G3481gat);
nor NOR2_1299 (G3664gat, G3556gat, G3608gat);
nor NOR2_1300 (G3665gat, G3608gat, G3486gat);
nor NOR2_1301 (G3666gat, G3559gat, G3612gat);
nor NOR2_1302 (G3667gat, G3612gat, G3491gat);
nor NOR2_1303 (G3668gat, G3562gat, G3616gat);
nor NOR2_1304 (G3669gat, G3616gat, G3496gat);
nor NOR2_1305 (G3670gat, G3565gat, G3620gat);
nor NOR2_1306 (G3671gat, G3620gat, G3501gat);
nor NOR2_1307 (G3672gat, G3568gat, G3624gat);
nor NOR2_1308 (G3673gat, G3624gat, G3506gat);
nor NOR2_1309 (G3674gat, G3571gat, G3628gat);
nor NOR2_1310 (G3675gat, G3628gat, G3511gat);
nor NOR2_1311 (G3676gat, G3574gat, G3632gat);
nor NOR2_1312 (G3677gat, G3632gat, G3516gat);
nor NOR2_1313 (G3678gat, G3636gat, G3637gat);
nor NOR2_1314 (G3681gat, G3638gat, G999gat);
nor NOR2_1315 (G3685gat, G3583gat, G3641gat);
nor NOR2_1316 (G3686gat, G3641gat, G1047gat);
nor NOR2_1317 (G3687gat, G3461gat, G3641gat);
nor NOR2_1318 (G3690gat, G3645gat, G3646gat);
nor NOR2_1319 (G3693gat, G3650gat, G3647gat);
nor NOR2_1320 (G3697gat, G3595gat, G3653gat);
nor NOR2_1321 (G3698gat, G3653gat, G3592gat);
nor NOR2_1322 (G3699gat, G3657gat, G3658gat);
nor NOR2_1323 (G3702gat, G3659gat, G1242gat);
nor NOR2_1324 (G3706gat, G3662gat, G3663gat);
nor NOR2_1325 (G3709gat, G3664gat, G3665gat);
nor NOR2_1326 (G3712gat, G3666gat, G3667gat);
nor NOR2_1327 (G3715gat, G3668gat, G3669gat);
nor NOR2_1328 (G3718gat, G3670gat, G3671gat);
nor NOR2_1329 (G3721gat, G3672gat, G3673gat);
nor NOR2_1330 (G3724gat, G3674gat, G3675gat);
nor NOR2_1331 (G3727gat, G3676gat, G3677gat);
nor NOR2_1332 (G3730gat, G3678gat, G951gat);
nor NOR2_1333 (G3734gat, G3638gat, G3681gat);
nor NOR2_1334 (G3735gat, G3681gat, G999gat);
nor NOR2_1335 (G3736gat, G3527gat, G3681gat);
nor NOR2_1336 (G3739gat, G3685gat, G3686gat);
nor NOR2_1337 (G3742gat, G3690gat, G3687gat);
nor NOR2_1338 (G3746gat, G3650gat, G3693gat);
nor NOR2_1339 (G3747gat, G3693gat, G3647gat);
nor NOR2_1340 (G3748gat, G3697gat, G3698gat);
nor NOR2_1341 (G3751gat, G3699gat, G1194gat);
nor NOR2_1342 (G3755gat, G3659gat, G3702gat);
nor NOR2_1343 (G3756gat, G3702gat, G1242gat);
nor NOR2_1344 (G3757gat, G3548gat, G3702gat);
nor NOR2_1345 (G3760gat, G3706gat, G567gat);
nor NOR2_1346 (G3764gat, G3709gat, G615gat);
nor NOR2_1347 (G3768gat, G3712gat, G663gat);
nor NOR2_1348 (G3772gat, G3715gat, G711gat);
nor NOR2_1349 (G3776gat, G3718gat, G759gat);
nor NOR2_1350 (G3780gat, G3721gat, G807gat);
nor NOR2_1351 (G3784gat, G3724gat, G855gat);
nor NOR2_1352 (G3788gat, G3727gat, G903gat);
nor NOR2_1353 (G3792gat, G3678gat, G3730gat);
nor NOR2_1354 (G3793gat, G3730gat, G951gat);
nor NOR2_1355 (G3794gat, G3577gat, G3730gat);
nor NOR2_1356 (G3797gat, G3734gat, G3735gat);
nor NOR2_1357 (G3800gat, G3739gat, G3736gat);
nor NOR2_1358 (G3804gat, G3690gat, G3742gat);
nor NOR2_1359 (G3805gat, G3742gat, G3687gat);
nor NOR2_1360 (G3806gat, G3746gat, G3747gat);
nor NOR2_1361 (G3809gat, G3748gat, G1146gat);
nor NOR2_1362 (G3813gat, G3699gat, G3751gat);
nor NOR2_1363 (G3814gat, G3751gat, G1194gat);
nor NOR2_1364 (G3815gat, G3598gat, G3751gat);
nor NOR2_1365 (G3818gat, G3755gat, G3756gat);
nor NOR2_1366 (G3821gat, G1290gat, G3757gat);
nor NOR2_1367 (G3825gat, G3706gat, G3760gat);
nor NOR2_1368 (G3826gat, G3760gat, G567gat);
nor NOR2_1369 (G3827gat, G3604gat, G3760gat);
nor NOR2_1370 (G3830gat, G3709gat, G3764gat);
nor NOR2_1371 (G3831gat, G3764gat, G615gat);
nor NOR2_1372 (G3832gat, G3608gat, G3764gat);
nor NOR2_1373 (G3835gat, G3712gat, G3768gat);
nor NOR2_1374 (G3836gat, G3768gat, G663gat);
nor NOR2_1375 (G3837gat, G3612gat, G3768gat);
nor NOR2_1376 (G3840gat, G3715gat, G3772gat);
nor NOR2_1377 (G3841gat, G3772gat, G711gat);
nor NOR2_1378 (G3842gat, G3616gat, G3772gat);
nor NOR2_1379 (G3845gat, G3718gat, G3776gat);
nor NOR2_1380 (G3846gat, G3776gat, G759gat);
nor NOR2_1381 (G3847gat, G3620gat, G3776gat);
nor NOR2_1382 (G3850gat, G3721gat, G3780gat);
nor NOR2_1383 (G3851gat, G3780gat, G807gat);
nor NOR2_1384 (G3852gat, G3624gat, G3780gat);
nor NOR2_1385 (G3855gat, G3724gat, G3784gat);
nor NOR2_1386 (G3856gat, G3784gat, G855gat);
nor NOR2_1387 (G3857gat, G3628gat, G3784gat);
nor NOR2_1388 (G3860gat, G3727gat, G3788gat);
nor NOR2_1389 (G3861gat, G3788gat, G903gat);
nor NOR2_1390 (G3862gat, G3632gat, G3788gat);
nor NOR2_1391 (G3865gat, G3792gat, G3793gat);
nor NOR2_1392 (G3868gat, G3797gat, G3794gat);
nor NOR2_1393 (G3872gat, G3739gat, G3800gat);
nor NOR2_1394 (G3873gat, G3800gat, G3736gat);
nor NOR2_1395 (G3874gat, G3804gat, G3805gat);
nor NOR2_1396 (G3877gat, G3806gat, G1098gat);
nor NOR2_1397 (G3881gat, G3748gat, G3809gat);
nor NOR2_1398 (G3882gat, G3809gat, G1146gat);
nor NOR2_1399 (G3883gat, G3653gat, G3809gat);
nor NOR2_1400 (G3886gat, G3813gat, G3814gat);
nor NOR2_1401 (G3889gat, G3818gat, G3815gat);
nor NOR2_1402 (G3893gat, G1290gat, G3821gat);
nor NOR2_1403 (G3894gat, G3821gat, G3757gat);
nor NOR2_1404 (G3895gat, G3825gat, G3826gat);
nor NOR2_1405 (G3896gat, G3830gat, G3831gat);
nor NOR2_1406 (G3899gat, G3835gat, G3836gat);
nor NOR2_1407 (G3902gat, G3840gat, G3841gat);
nor NOR2_1408 (G3905gat, G3845gat, G3846gat);
nor NOR2_1409 (G3908gat, G3850gat, G3851gat);
nor NOR2_1410 (G3911gat, G3855gat, G3856gat);
nor NOR2_1411 (G3914gat, G3860gat, G3861gat);
nor NOR2_1412 (G3917gat, G3865gat, G3862gat);
nor NOR2_1413 (G3921gat, G3797gat, G3868gat);
nor NOR2_1414 (G3922gat, G3868gat, G3794gat);
nor NOR2_1415 (G3923gat, G3872gat, G3873gat);
nor NOR2_1416 (G3926gat, G3874gat, G1050gat);
nor NOR2_1417 (G3930gat, G3806gat, G3877gat);
nor NOR2_1418 (G3931gat, G3877gat, G1098gat);
nor NOR2_1419 (G3932gat, G3693gat, G3877gat);
nor NOR2_1420 (G3935gat, G3881gat, G3882gat);
nor NOR2_1421 (G3938gat, G3886gat, G3883gat);
nor NOR2_1422 (G3942gat, G3818gat, G3889gat);
nor NOR2_1423 (G3943gat, G3889gat, G3815gat);
nor NOR2_1424 (G3944gat, G3893gat, G3894gat);
nor NOR2_1425 (G3947gat, G3896gat, G3827gat);
nor NOR2_1426 (G3951gat, G3899gat, G3832gat);
nor NOR2_1427 (G3955gat, G3902gat, G3837gat);
nor NOR2_1428 (G3959gat, G3905gat, G3842gat);
nor NOR2_1429 (G3963gat, G3908gat, G3847gat);
nor NOR2_1430 (G3967gat, G3911gat, G3852gat);
nor NOR2_1431 (G3971gat, G3914gat, G3857gat);
nor NOR2_1432 (G3975gat, G3865gat, G3917gat);
nor NOR2_1433 (G3976gat, G3917gat, G3862gat);
nor NOR2_1434 (G3977gat, G3921gat, G3922gat);
nor NOR2_1435 (G3980gat, G3923gat, G1002gat);
nor NOR2_1436 (G3984gat, G3874gat, G3926gat);
nor NOR2_1437 (G3985gat, G3926gat, G1050gat);
nor NOR2_1438 (G3986gat, G3742gat, G3926gat);
nor NOR2_1439 (G3989gat, G3930gat, G3931gat);
nor NOR2_1440 (G3992gat, G3935gat, G3932gat);
nor NOR2_1441 (G3996gat, G3886gat, G3938gat);
nor NOR2_1442 (G3997gat, G3938gat, G3883gat);
nor NOR2_1443 (G3998gat, G3942gat, G3943gat);
nor NOR2_1444 (G4001gat, G3944gat, G1245gat);
nor NOR2_1445 (G4005gat, G3896gat, G3947gat);
nor NOR2_1446 (G4006gat, G3947gat, G3827gat);
nor NOR2_1447 (G4007gat, G3899gat, G3951gat);
nor NOR2_1448 (G4008gat, G3951gat, G3832gat);
nor NOR2_1449 (G4009gat, G3902gat, G3955gat);
nor NOR2_1450 (G4010gat, G3955gat, G3837gat);
nor NOR2_1451 (G4011gat, G3905gat, G3959gat);
nor NOR2_1452 (G4012gat, G3959gat, G3842gat);
nor NOR2_1453 (G4013gat, G3908gat, G3963gat);
nor NOR2_1454 (G4014gat, G3963gat, G3847gat);
nor NOR2_1455 (G4015gat, G3911gat, G3967gat);
nor NOR2_1456 (G4016gat, G3967gat, G3852gat);
nor NOR2_1457 (G4017gat, G3914gat, G3971gat);
nor NOR2_1458 (G4018gat, G3971gat, G3857gat);
nor NOR2_1459 (G4019gat, G3975gat, G3976gat);
nor NOR2_1460 (G4022gat, G3977gat, G954gat);
nor NOR2_1461 (G4026gat, G3923gat, G3980gat);
nor NOR2_1462 (G4027gat, G3980gat, G1002gat);
nor NOR2_1463 (G4028gat, G3800gat, G3980gat);
nor NOR2_1464 (G4031gat, G3984gat, G3985gat);
nor NOR2_1465 (G4034gat, G3989gat, G3986gat);
nor NOR2_1466 (G4038gat, G3935gat, G3992gat);
nor NOR2_1467 (G4039gat, G3992gat, G3932gat);
nor NOR2_1468 (G4040gat, G3996gat, G3997gat);
nor NOR2_1469 (G4043gat, G3998gat, G1197gat);
nor NOR2_1470 (G4047gat, G3944gat, G4001gat);
nor NOR2_1471 (G4048gat, G4001gat, G1245gat);
nor NOR2_1472 (G4049gat, G3821gat, G4001gat);
nor NOR2_1473 (G4052gat, G4005gat, G4006gat);
nor NOR2_1474 (G4055gat, G4007gat, G4008gat);
nor NOR2_1475 (G4058gat, G4009gat, G4010gat);
nor NOR2_1476 (G4061gat, G4011gat, G4012gat);
nor NOR2_1477 (G4064gat, G4013gat, G4014gat);
nor NOR2_1478 (G4067gat, G4015gat, G4016gat);
nor NOR2_1479 (G4070gat, G4017gat, G4018gat);
nor NOR2_1480 (G4073gat, G4019gat, G906gat);
nor NOR2_1481 (G4077gat, G3977gat, G4022gat);
nor NOR2_1482 (G4078gat, G4022gat, G954gat);
nor NOR2_1483 (G4079gat, G3868gat, G4022gat);
nor NOR2_1484 (G4082gat, G4026gat, G4027gat);
nor NOR2_1485 (G4085gat, G4031gat, G4028gat);
nor NOR2_1486 (G4089gat, G3989gat, G4034gat);
nor NOR2_1487 (G4090gat, G4034gat, G3986gat);
nor NOR2_1488 (G4091gat, G4038gat, G4039gat);
nor NOR2_1489 (G4094gat, G4040gat, G1149gat);
nor NOR2_1490 (G4098gat, G3998gat, G4043gat);
nor NOR2_1491 (G4099gat, G4043gat, G1197gat);
nor NOR2_1492 (G4100gat, G3889gat, G4043gat);
nor NOR2_1493 (G4103gat, G4047gat, G4048gat);
nor NOR2_1494 (G4106gat, G1293gat, G4049gat);
nor NOR2_1495 (G4110gat, G4052gat, G570gat);
nor NOR2_1496 (G4114gat, G4055gat, G618gat);
nor NOR2_1497 (G4118gat, G4058gat, G666gat);
nor NOR2_1498 (G4122gat, G4061gat, G714gat);
nor NOR2_1499 (G4126gat, G4064gat, G762gat);
nor NOR2_1500 (G4130gat, G4067gat, G810gat);
nor NOR2_1501 (G4134gat, G4070gat, G858gat);
nor NOR2_1502 (G4138gat, G4019gat, G4073gat);
nor NOR2_1503 (G4139gat, G4073gat, G906gat);
nor NOR2_1504 (G4140gat, G3917gat, G4073gat);
nor NOR2_1505 (G4143gat, G4077gat, G4078gat);
nor NOR2_1506 (G4146gat, G4082gat, G4079gat);
nor NOR2_1507 (G4150gat, G4031gat, G4085gat);
nor NOR2_1508 (G4151gat, G4085gat, G4028gat);
nor NOR2_1509 (G4152gat, G4089gat, G4090gat);
nor NOR2_1510 (G4155gat, G4091gat, G1101gat);
nor NOR2_1511 (G4159gat, G4040gat, G4094gat);
nor NOR2_1512 (G4160gat, G4094gat, G1149gat);
nor NOR2_1513 (G4161gat, G3938gat, G4094gat);
nor NOR2_1514 (G4164gat, G4098gat, G4099gat);
nor NOR2_1515 (G4167gat, G4103gat, G4100gat);
nor NOR2_1516 (G4171gat, G1293gat, G4106gat);
nor NOR2_1517 (G4172gat, G4106gat, G4049gat);
nor NOR2_1518 (G4173gat, G4052gat, G4110gat);
nor NOR2_1519 (G4174gat, G4110gat, G570gat);
nor NOR2_1520 (G4175gat, G3947gat, G4110gat);
nor NOR2_1521 (G4178gat, G4055gat, G4114gat);
nor NOR2_1522 (G4179gat, G4114gat, G618gat);
nor NOR2_1523 (G4180gat, G3951gat, G4114gat);
nor NOR2_1524 (G4183gat, G4058gat, G4118gat);
nor NOR2_1525 (G4184gat, G4118gat, G666gat);
nor NOR2_1526 (G4185gat, G3955gat, G4118gat);
nor NOR2_1527 (G4188gat, G4061gat, G4122gat);
nor NOR2_1528 (G4189gat, G4122gat, G714gat);
nor NOR2_1529 (G4190gat, G3959gat, G4122gat);
nor NOR2_1530 (G4193gat, G4064gat, G4126gat);
nor NOR2_1531 (G4194gat, G4126gat, G762gat);
nor NOR2_1532 (G4195gat, G3963gat, G4126gat);
nor NOR2_1533 (G4198gat, G4067gat, G4130gat);
nor NOR2_1534 (G4199gat, G4130gat, G810gat);
nor NOR2_1535 (G4200gat, G3967gat, G4130gat);
nor NOR2_1536 (G4203gat, G4070gat, G4134gat);
nor NOR2_1537 (G4204gat, G4134gat, G858gat);
nor NOR2_1538 (G4205gat, G3971gat, G4134gat);
nor NOR2_1539 (G4208gat, G4138gat, G4139gat);
nor NOR2_1540 (G4211gat, G4143gat, G4140gat);
nor NOR2_1541 (G4215gat, G4082gat, G4146gat);
nor NOR2_1542 (G4216gat, G4146gat, G4079gat);
nor NOR2_1543 (G4217gat, G4150gat, G4151gat);
nor NOR2_1544 (G4220gat, G4152gat, G1053gat);
nor NOR2_1545 (G4224gat, G4091gat, G4155gat);
nor NOR2_1546 (G4225gat, G4155gat, G1101gat);
nor NOR2_1547 (G4226gat, G3992gat, G4155gat);
nor NOR2_1548 (G4229gat, G4159gat, G4160gat);
nor NOR2_1549 (G4232gat, G4164gat, G4161gat);
nor NOR2_1550 (G4236gat, G4103gat, G4167gat);
nor NOR2_1551 (G4237gat, G4167gat, G4100gat);
nor NOR2_1552 (G4238gat, G4171gat, G4172gat);
nor NOR2_1553 (G4241gat, G4173gat, G4174gat);
nor NOR2_1554 (G4242gat, G4178gat, G4179gat);
nor NOR2_1555 (G4245gat, G4183gat, G4184gat);
nor NOR2_1556 (G4248gat, G4188gat, G4189gat);
nor NOR2_1557 (G4251gat, G4193gat, G4194gat);
nor NOR2_1558 (G4254gat, G4198gat, G4199gat);
nor NOR2_1559 (G4257gat, G4203gat, G4204gat);
nor NOR2_1560 (G4260gat, G4208gat, G4205gat);
nor NOR2_1561 (G4264gat, G4143gat, G4211gat);
nor NOR2_1562 (G4265gat, G4211gat, G4140gat);
nor NOR2_1563 (G4266gat, G4215gat, G4216gat);
nor NOR2_1564 (G4269gat, G4217gat, G1005gat);
nor NOR2_1565 (G4273gat, G4152gat, G4220gat);
nor NOR2_1566 (G4274gat, G4220gat, G1053gat);
nor NOR2_1567 (G4275gat, G4034gat, G4220gat);
nor NOR2_1568 (G4278gat, G4224gat, G4225gat);
nor NOR2_1569 (G4281gat, G4229gat, G4226gat);
nor NOR2_1570 (G4285gat, G4164gat, G4232gat);
nor NOR2_1571 (G4286gat, G4232gat, G4161gat);
nor NOR2_1572 (G4287gat, G4236gat, G4237gat);
nor NOR2_1573 (G4290gat, G4238gat, G1248gat);
nor NOR2_1574 (G4294gat, G4242gat, G4175gat);
nor NOR2_1575 (G4298gat, G4245gat, G4180gat);
nor NOR2_1576 (G4302gat, G4248gat, G4185gat);
nor NOR2_1577 (G4306gat, G4251gat, G4190gat);
nor NOR2_1578 (G4310gat, G4254gat, G4195gat);
nor NOR2_1579 (G4314gat, G4257gat, G4200gat);
nor NOR2_1580 (G4318gat, G4208gat, G4260gat);
nor NOR2_1581 (G4319gat, G4260gat, G4205gat);
nor NOR2_1582 (G4320gat, G4264gat, G4265gat);
nor NOR2_1583 (G4323gat, G4266gat, G957gat);
nor NOR2_1584 (G4327gat, G4217gat, G4269gat);
nor NOR2_1585 (G4328gat, G4269gat, G1005gat);
nor NOR2_1586 (G4329gat, G4085gat, G4269gat);
nor NOR2_1587 (G4332gat, G4273gat, G4274gat);
nor NOR2_1588 (G4335gat, G4278gat, G4275gat);
nor NOR2_1589 (G4339gat, G4229gat, G4281gat);
nor NOR2_1590 (G4340gat, G4281gat, G4226gat);
nor NOR2_1591 (G4341gat, G4285gat, G4286gat);
nor NOR2_1592 (G4344gat, G4287gat, G1200gat);
nor NOR2_1593 (G4348gat, G4238gat, G4290gat);
nor NOR2_1594 (G4349gat, G4290gat, G1248gat);
nor NOR2_1595 (G4350gat, G4106gat, G4290gat);
nor NOR2_1596 (G4353gat, G4242gat, G4294gat);
nor NOR2_1597 (G4354gat, G4294gat, G4175gat);
nor NOR2_1598 (G4355gat, G4245gat, G4298gat);
nor NOR2_1599 (G4356gat, G4298gat, G4180gat);
nor NOR2_1600 (G4357gat, G4248gat, G4302gat);
nor NOR2_1601 (G4358gat, G4302gat, G4185gat);
nor NOR2_1602 (G4359gat, G4251gat, G4306gat);
nor NOR2_1603 (G4360gat, G4306gat, G4190gat);
nor NOR2_1604 (G4361gat, G4254gat, G4310gat);
nor NOR2_1605 (G4362gat, G4310gat, G4195gat);
nor NOR2_1606 (G4363gat, G4257gat, G4314gat);
nor NOR2_1607 (G4364gat, G4314gat, G4200gat);
nor NOR2_1608 (G4365gat, G4318gat, G4319gat);
nor NOR2_1609 (G4368gat, G4320gat, G909gat);
nor NOR2_1610 (G4372gat, G4266gat, G4323gat);
nor NOR2_1611 (G4373gat, G4323gat, G957gat);
nor NOR2_1612 (G4374gat, G4146gat, G4323gat);
nor NOR2_1613 (G4377gat, G4327gat, G4328gat);
nor NOR2_1614 (G4380gat, G4332gat, G4329gat);
nor NOR2_1615 (G4384gat, G4278gat, G4335gat);
nor NOR2_1616 (G4385gat, G4335gat, G4275gat);
nor NOR2_1617 (G4386gat, G4339gat, G4340gat);
nor NOR2_1618 (G4389gat, G4341gat, G1152gat);
nor NOR2_1619 (G4393gat, G4287gat, G4344gat);
nor NOR2_1620 (G4394gat, G4344gat, G1200gat);
nor NOR2_1621 (G4395gat, G4167gat, G4344gat);
nor NOR2_1622 (G4398gat, G4348gat, G4349gat);
nor NOR2_1623 (G4401gat, G1296gat, G4350gat);
nor NOR2_1624 (G4405gat, G4353gat, G4354gat);
nor NOR2_1625 (G4408gat, G4355gat, G4356gat);
nor NOR2_1626 (G4411gat, G4357gat, G4358gat);
nor NOR2_1627 (G4414gat, G4359gat, G4360gat);
nor NOR2_1628 (G4417gat, G4361gat, G4362gat);
nor NOR2_1629 (G4420gat, G4363gat, G4364gat);
nor NOR2_1630 (G4423gat, G4365gat, G861gat);
nor NOR2_1631 (G4427gat, G4320gat, G4368gat);
nor NOR2_1632 (G4428gat, G4368gat, G909gat);
nor NOR2_1633 (G4429gat, G4211gat, G4368gat);
nor NOR2_1634 (G4432gat, G4372gat, G4373gat);
nor NOR2_1635 (G4435gat, G4377gat, G4374gat);
nor NOR2_1636 (G4439gat, G4332gat, G4380gat);
nor NOR2_1637 (G4440gat, G4380gat, G4329gat);
nor NOR2_1638 (G4441gat, G4384gat, G4385gat);
nor NOR2_1639 (G4444gat, G4386gat, G1104gat);
nor NOR2_1640 (G4448gat, G4341gat, G4389gat);
nor NOR2_1641 (G4449gat, G4389gat, G1152gat);
nor NOR2_1642 (G4450gat, G4232gat, G4389gat);
nor NOR2_1643 (G4453gat, G4393gat, G4394gat);
nor NOR2_1644 (G4456gat, G4398gat, G4395gat);
nor NOR2_1645 (G4460gat, G1296gat, G4401gat);
nor NOR2_1646 (G4461gat, G4401gat, G4350gat);
nor NOR2_1647 (G4462gat, G4405gat, G573gat);
nor NOR2_1648 (G4466gat, G4408gat, G621gat);
nor NOR2_1649 (G4470gat, G4411gat, G669gat);
nor NOR2_1650 (G4474gat, G4414gat, G717gat);
nor NOR2_1651 (G4478gat, G4417gat, G765gat);
nor NOR2_1652 (G4482gat, G4420gat, G813gat);
nor NOR2_1653 (G4486gat, G4365gat, G4423gat);
nor NOR2_1654 (G4487gat, G4423gat, G861gat);
nor NOR2_1655 (G4488gat, G4260gat, G4423gat);
nor NOR2_1656 (G4491gat, G4427gat, G4428gat);
nor NOR2_1657 (G4494gat, G4432gat, G4429gat);
nor NOR2_1658 (G4498gat, G4377gat, G4435gat);
nor NOR2_1659 (G4499gat, G4435gat, G4374gat);
nor NOR2_1660 (G4500gat, G4439gat, G4440gat);
nor NOR2_1661 (G4503gat, G4441gat, G1056gat);
nor NOR2_1662 (G4507gat, G4386gat, G4444gat);
nor NOR2_1663 (G4508gat, G4444gat, G1104gat);
nor NOR2_1664 (G4509gat, G4281gat, G4444gat);
nor NOR2_1665 (G4512gat, G4448gat, G4449gat);
nor NOR2_1666 (G4515gat, G4453gat, G4450gat);
nor NOR2_1667 (G4519gat, G4398gat, G4456gat);
nor NOR2_1668 (G4520gat, G4456gat, G4395gat);
nor NOR2_1669 (G4521gat, G4460gat, G4461gat);
nor NOR2_1670 (G4524gat, G4405gat, G4462gat);
nor NOR2_1671 (G4525gat, G4462gat, G573gat);
nor NOR2_1672 (G4526gat, G4294gat, G4462gat);
nor NOR2_1673 (G4529gat, G4408gat, G4466gat);
nor NOR2_1674 (G4530gat, G4466gat, G621gat);
nor NOR2_1675 (G4531gat, G4298gat, G4466gat);
nor NOR2_1676 (G4534gat, G4411gat, G4470gat);
nor NOR2_1677 (G4535gat, G4470gat, G669gat);
nor NOR2_1678 (G4536gat, G4302gat, G4470gat);
nor NOR2_1679 (G4539gat, G4414gat, G4474gat);
nor NOR2_1680 (G4540gat, G4474gat, G717gat);
nor NOR2_1681 (G4541gat, G4306gat, G4474gat);
nor NOR2_1682 (G4544gat, G4417gat, G4478gat);
nor NOR2_1683 (G4545gat, G4478gat, G765gat);
nor NOR2_1684 (G4546gat, G4310gat, G4478gat);
nor NOR2_1685 (G4549gat, G4420gat, G4482gat);
nor NOR2_1686 (G4550gat, G4482gat, G813gat);
nor NOR2_1687 (G4551gat, G4314gat, G4482gat);
nor NOR2_1688 (G4554gat, G4486gat, G4487gat);
nor NOR2_1689 (G4557gat, G4491gat, G4488gat);
nor NOR2_1690 (G4561gat, G4432gat, G4494gat);
nor NOR2_1691 (G4562gat, G4494gat, G4429gat);
nor NOR2_1692 (G4563gat, G4498gat, G4499gat);
nor NOR2_1693 (G4566gat, G4500gat, G1008gat);
nor NOR2_1694 (G4570gat, G4441gat, G4503gat);
nor NOR2_1695 (G4571gat, G4503gat, G1056gat);
nor NOR2_1696 (G4572gat, G4335gat, G4503gat);
nor NOR2_1697 (G4575gat, G4507gat, G4508gat);
nor NOR2_1698 (G4578gat, G4512gat, G4509gat);
nor NOR2_1699 (G4582gat, G4453gat, G4515gat);
nor NOR2_1700 (G4583gat, G4515gat, G4450gat);
nor NOR2_1701 (G4584gat, G4519gat, G4520gat);
nor NOR2_1702 (G4587gat, G4521gat, G1251gat);
nor NOR2_1703 (G4591gat, G4524gat, G4525gat);
nor NOR2_1704 (G4592gat, G4529gat, G4530gat);
nor NOR2_1705 (G4595gat, G4534gat, G4535gat);
nor NOR2_1706 (G4598gat, G4539gat, G4540gat);
nor NOR2_1707 (G4601gat, G4544gat, G4545gat);
nor NOR2_1708 (G4604gat, G4549gat, G4550gat);
nor NOR2_1709 (G4607gat, G4554gat, G4551gat);
nor NOR2_1710 (G4611gat, G4491gat, G4557gat);
nor NOR2_1711 (G4612gat, G4557gat, G4488gat);
nor NOR2_1712 (G4613gat, G4561gat, G4562gat);
nor NOR2_1713 (G4616gat, G4563gat, G960gat);
nor NOR2_1714 (G4620gat, G4500gat, G4566gat);
nor NOR2_1715 (G4621gat, G4566gat, G1008gat);
nor NOR2_1716 (G4622gat, G4380gat, G4566gat);
nor NOR2_1717 (G4625gat, G4570gat, G4571gat);
nor NOR2_1718 (G4628gat, G4575gat, G4572gat);
nor NOR2_1719 (G4632gat, G4512gat, G4578gat);
nor NOR2_1720 (G4633gat, G4578gat, G4509gat);
nor NOR2_1721 (G4634gat, G4582gat, G4583gat);
nor NOR2_1722 (G4637gat, G4584gat, G1203gat);
nor NOR2_1723 (G4641gat, G4521gat, G4587gat);
nor NOR2_1724 (G4642gat, G4587gat, G1251gat);
nor NOR2_1725 (G4643gat, G4401gat, G4587gat);
nor NOR2_1726 (G4646gat, G4592gat, G4526gat);
nor NOR2_1727 (G4650gat, G4595gat, G4531gat);
nor NOR2_1728 (G4654gat, G4598gat, G4536gat);
nor NOR2_1729 (G4658gat, G4601gat, G4541gat);
nor NOR2_1730 (G4662gat, G4604gat, G4546gat);
nor NOR2_1731 (G4666gat, G4554gat, G4607gat);
nor NOR2_1732 (G4667gat, G4607gat, G4551gat);
nor NOR2_1733 (G4668gat, G4611gat, G4612gat);
nor NOR2_1734 (G4671gat, G4613gat, G912gat);
nor NOR2_1735 (G4675gat, G4563gat, G4616gat);
nor NOR2_1736 (G4676gat, G4616gat, G960gat);
nor NOR2_1737 (G4677gat, G4435gat, G4616gat);
nor NOR2_1738 (G4680gat, G4620gat, G4621gat);
nor NOR2_1739 (G4683gat, G4625gat, G4622gat);
nor NOR2_1740 (G4687gat, G4575gat, G4628gat);
nor NOR2_1741 (G4688gat, G4628gat, G4572gat);
nor NOR2_1742 (G4689gat, G4632gat, G4633gat);
nor NOR2_1743 (G4692gat, G4634gat, G1155gat);
nor NOR2_1744 (G4696gat, G4584gat, G4637gat);
nor NOR2_1745 (G4697gat, G4637gat, G1203gat);
nor NOR2_1746 (G4698gat, G4456gat, G4637gat);
nor NOR2_1747 (G4701gat, G4641gat, G4642gat);
nor NOR2_1748 (G4704gat, G1299gat, G4643gat);
nor NOR2_1749 (G4708gat, G4592gat, G4646gat);
nor NOR2_1750 (G4709gat, G4646gat, G4526gat);
nor NOR2_1751 (G4710gat, G4595gat, G4650gat);
nor NOR2_1752 (G4711gat, G4650gat, G4531gat);
nor NOR2_1753 (G4712gat, G4598gat, G4654gat);
nor NOR2_1754 (G4713gat, G4654gat, G4536gat);
nor NOR2_1755 (G4714gat, G4601gat, G4658gat);
nor NOR2_1756 (G4715gat, G4658gat, G4541gat);
nor NOR2_1757 (G4716gat, G4604gat, G4662gat);
nor NOR2_1758 (G4717gat, G4662gat, G4546gat);
nor NOR2_1759 (G4718gat, G4666gat, G4667gat);
nor NOR2_1760 (G4721gat, G4668gat, G864gat);
nor NOR2_1761 (G4725gat, G4613gat, G4671gat);
nor NOR2_1762 (G4726gat, G4671gat, G912gat);
nor NOR2_1763 (G4727gat, G4494gat, G4671gat);
nor NOR2_1764 (G4730gat, G4675gat, G4676gat);
nor NOR2_1765 (G4733gat, G4680gat, G4677gat);
nor NOR2_1766 (G4737gat, G4625gat, G4683gat);
nor NOR2_1767 (G4738gat, G4683gat, G4622gat);
nor NOR2_1768 (G4739gat, G4687gat, G4688gat);
nor NOR2_1769 (G4742gat, G4689gat, G1107gat);
nor NOR2_1770 (G4746gat, G4634gat, G4692gat);
nor NOR2_1771 (G4747gat, G4692gat, G1155gat);
nor NOR2_1772 (G4748gat, G4515gat, G4692gat);
nor NOR2_1773 (G4751gat, G4696gat, G4697gat);
nor NOR2_1774 (G4754gat, G4701gat, G4698gat);
nor NOR2_1775 (G4758gat, G1299gat, G4704gat);
nor NOR2_1776 (G4759gat, G4704gat, G4643gat);
nor NOR2_1777 (G4760gat, G4708gat, G4709gat);
nor NOR2_1778 (G4763gat, G4710gat, G4711gat);
nor NOR2_1779 (G4766gat, G4712gat, G4713gat);
nor NOR2_1780 (G4769gat, G4714gat, G4715gat);
nor NOR2_1781 (G4772gat, G4716gat, G4717gat);
nor NOR2_1782 (G4775gat, G4718gat, G816gat);
nor NOR2_1783 (G4779gat, G4668gat, G4721gat);
nor NOR2_1784 (G4780gat, G4721gat, G864gat);
nor NOR2_1785 (G4781gat, G4557gat, G4721gat);
nor NOR2_1786 (G4784gat, G4725gat, G4726gat);
nor NOR2_1787 (G4787gat, G4730gat, G4727gat);
nor NOR2_1788 (G4791gat, G4680gat, G4733gat);
nor NOR2_1789 (G4792gat, G4733gat, G4677gat);
nor NOR2_1790 (G4793gat, G4737gat, G4738gat);
nor NOR2_1791 (G4796gat, G4739gat, G1059gat);
nor NOR2_1792 (G4800gat, G4689gat, G4742gat);
nor NOR2_1793 (G4801gat, G4742gat, G1107gat);
nor NOR2_1794 (G4802gat, G4578gat, G4742gat);
nor NOR2_1795 (G4805gat, G4746gat, G4747gat);
nor NOR2_1796 (G4808gat, G4751gat, G4748gat);
nor NOR2_1797 (G4812gat, G4701gat, G4754gat);
nor NOR2_1798 (G4813gat, G4754gat, G4698gat);
nor NOR2_1799 (G4814gat, G4758gat, G4759gat);
nor NOR2_1800 (G4817gat, G4760gat, G576gat);
nor NOR2_1801 (G4821gat, G4763gat, G624gat);
nor NOR2_1802 (G4825gat, G4766gat, G672gat);
nor NOR2_1803 (G4829gat, G4769gat, G720gat);
nor NOR2_1804 (G4833gat, G4772gat, G768gat);
nor NOR2_1805 (G4837gat, G4718gat, G4775gat);
nor NOR2_1806 (G4838gat, G4775gat, G816gat);
nor NOR2_1807 (G4839gat, G4607gat, G4775gat);
nor NOR2_1808 (G4842gat, G4779gat, G4780gat);
nor NOR2_1809 (G4845gat, G4784gat, G4781gat);
nor NOR2_1810 (G4849gat, G4730gat, G4787gat);
nor NOR2_1811 (G4850gat, G4787gat, G4727gat);
nor NOR2_1812 (G4851gat, G4791gat, G4792gat);
nor NOR2_1813 (G4854gat, G4793gat, G1011gat);
nor NOR2_1814 (G4858gat, G4739gat, G4796gat);
nor NOR2_1815 (G4859gat, G4796gat, G1059gat);
nor NOR2_1816 (G4860gat, G4628gat, G4796gat);
nor NOR2_1817 (G4863gat, G4800gat, G4801gat);
nor NOR2_1818 (G4866gat, G4805gat, G4802gat);
nor NOR2_1819 (G4870gat, G4751gat, G4808gat);
nor NOR2_1820 (G4871gat, G4808gat, G4748gat);
nor NOR2_1821 (G4872gat, G4812gat, G4813gat);
nor NOR2_1822 (G4875gat, G4814gat, G1254gat);
nor NOR2_1823 (G4879gat, G4760gat, G4817gat);
nor NOR2_1824 (G4880gat, G4817gat, G576gat);
nor NOR2_1825 (G4881gat, G4646gat, G4817gat);
nor NOR2_1826 (G4884gat, G4763gat, G4821gat);
nor NOR2_1827 (G4885gat, G4821gat, G624gat);
nor NOR2_1828 (G4886gat, G4650gat, G4821gat);
nor NOR2_1829 (G4889gat, G4766gat, G4825gat);
nor NOR2_1830 (G4890gat, G4825gat, G672gat);
nor NOR2_1831 (G4891gat, G4654gat, G4825gat);
nor NOR2_1832 (G4894gat, G4769gat, G4829gat);
nor NOR2_1833 (G4895gat, G4829gat, G720gat);
nor NOR2_1834 (G4896gat, G4658gat, G4829gat);
nor NOR2_1835 (G4899gat, G4772gat, G4833gat);
nor NOR2_1836 (G4900gat, G4833gat, G768gat);
nor NOR2_1837 (G4901gat, G4662gat, G4833gat);
nor NOR2_1838 (G4904gat, G4837gat, G4838gat);
nor NOR2_1839 (G4907gat, G4842gat, G4839gat);
nor NOR2_1840 (G4911gat, G4784gat, G4845gat);
nor NOR2_1841 (G4912gat, G4845gat, G4781gat);
nor NOR2_1842 (G4913gat, G4849gat, G4850gat);
nor NOR2_1843 (G4916gat, G4851gat, G963gat);
nor NOR2_1844 (G4920gat, G4793gat, G4854gat);
nor NOR2_1845 (G4921gat, G4854gat, G1011gat);
nor NOR2_1846 (G4922gat, G4683gat, G4854gat);
nor NOR2_1847 (G4925gat, G4858gat, G4859gat);
nor NOR2_1848 (G4928gat, G4863gat, G4860gat);
nor NOR2_1849 (G4932gat, G4805gat, G4866gat);
nor NOR2_1850 (G4933gat, G4866gat, G4802gat);
nor NOR2_1851 (G4934gat, G4870gat, G4871gat);
nor NOR2_1852 (G4937gat, G4872gat, G1206gat);
nor NOR2_1853 (G4941gat, G4814gat, G4875gat);
nor NOR2_1854 (G4942gat, G4875gat, G1254gat);
nor NOR2_1855 (G4943gat, G4704gat, G4875gat);
nor NOR2_1856 (G4946gat, G4879gat, G4880gat);
nor NOR2_1857 (G4947gat, G4884gat, G4885gat);
nor NOR2_1858 (G4950gat, G4889gat, G4890gat);
nor NOR2_1859 (G4953gat, G4894gat, G4895gat);
nor NOR2_1860 (G4956gat, G4899gat, G4900gat);
nor NOR2_1861 (G4959gat, G4904gat, G4901gat);
nor NOR2_1862 (G4963gat, G4842gat, G4907gat);
nor NOR2_1863 (G4964gat, G4907gat, G4839gat);
nor NOR2_1864 (G4965gat, G4911gat, G4912gat);
nor NOR2_1865 (G4968gat, G4913gat, G915gat);
nor NOR2_1866 (G4972gat, G4851gat, G4916gat);
nor NOR2_1867 (G4973gat, G4916gat, G963gat);
nor NOR2_1868 (G4974gat, G4733gat, G4916gat);
nor NOR2_1869 (G4977gat, G4920gat, G4921gat);
nor NOR2_1870 (G4980gat, G4925gat, G4922gat);
nor NOR2_1871 (G4984gat, G4863gat, G4928gat);
nor NOR2_1872 (G4985gat, G4928gat, G4860gat);
nor NOR2_1873 (G4986gat, G4932gat, G4933gat);
nor NOR2_1874 (G4989gat, G4934gat, G1158gat);
nor NOR2_1875 (G4993gat, G4872gat, G4937gat);
nor NOR2_1876 (G4994gat, G4937gat, G1206gat);
nor NOR2_1877 (G4995gat, G4754gat, G4937gat);
nor NOR2_1878 (G4998gat, G4941gat, G4942gat);
nor NOR2_1879 (G5001gat, G1302gat, G4943gat);
nor NOR2_1880 (G5005gat, G4947gat, G4881gat);
nor NOR2_1881 (G5009gat, G4950gat, G4886gat);
nor NOR2_1882 (G5013gat, G4953gat, G4891gat);
nor NOR2_1883 (G5017gat, G4956gat, G4896gat);
nor NOR2_1884 (G5021gat, G4904gat, G4959gat);
nor NOR2_1885 (G5022gat, G4959gat, G4901gat);
nor NOR2_1886 (G5023gat, G4963gat, G4964gat);
nor NOR2_1887 (G5026gat, G4965gat, G867gat);
nor NOR2_1888 (G5030gat, G4913gat, G4968gat);
nor NOR2_1889 (G5031gat, G4968gat, G915gat);
nor NOR2_1890 (G5032gat, G4787gat, G4968gat);
nor NOR2_1891 (G5035gat, G4972gat, G4973gat);
nor NOR2_1892 (G5038gat, G4977gat, G4974gat);
nor NOR2_1893 (G5042gat, G4925gat, G4980gat);
nor NOR2_1894 (G5043gat, G4980gat, G4922gat);
nor NOR2_1895 (G5044gat, G4984gat, G4985gat);
nor NOR2_1896 (G5047gat, G4986gat, G1110gat);
nor NOR2_1897 (G5051gat, G4934gat, G4989gat);
nor NOR2_1898 (G5052gat, G4989gat, G1158gat);
nor NOR2_1899 (G5053gat, G4808gat, G4989gat);
nor NOR2_1900 (G5056gat, G4993gat, G4994gat);
nor NOR2_1901 (G5059gat, G4998gat, G4995gat);
nor NOR2_1902 (G5063gat, G1302gat, G5001gat);
nor NOR2_1903 (G5064gat, G5001gat, G4943gat);
nor NOR2_1904 (G5065gat, G4947gat, G5005gat);
nor NOR2_1905 (G5066gat, G5005gat, G4881gat);
nor NOR2_1906 (G5067gat, G4950gat, G5009gat);
nor NOR2_1907 (G5068gat, G5009gat, G4886gat);
nor NOR2_1908 (G5069gat, G4953gat, G5013gat);
nor NOR2_1909 (G5070gat, G5013gat, G4891gat);
nor NOR2_1910 (G5071gat, G4956gat, G5017gat);
nor NOR2_1911 (G5072gat, G5017gat, G4896gat);
nor NOR2_1912 (G5073gat, G5021gat, G5022gat);
nor NOR2_1913 (G5076gat, G5023gat, G819gat);
nor NOR2_1914 (G5080gat, G4965gat, G5026gat);
nor NOR2_1915 (G5081gat, G5026gat, G867gat);
nor NOR2_1916 (G5082gat, G4845gat, G5026gat);
nor NOR2_1917 (G5085gat, G5030gat, G5031gat);
nor NOR2_1918 (G5088gat, G5035gat, G5032gat);
nor NOR2_1919 (G5092gat, G4977gat, G5038gat);
nor NOR2_1920 (G5093gat, G5038gat, G4974gat);
nor NOR2_1921 (G5094gat, G5042gat, G5043gat);
nor NOR2_1922 (G5097gat, G5044gat, G1062gat);
nor NOR2_1923 (G5101gat, G4986gat, G5047gat);
nor NOR2_1924 (G5102gat, G5047gat, G1110gat);
nor NOR2_1925 (G5103gat, G4866gat, G5047gat);
nor NOR2_1926 (G5106gat, G5051gat, G5052gat);
nor NOR2_1927 (G5109gat, G5056gat, G5053gat);
nor NOR2_1928 (G5113gat, G4998gat, G5059gat);
nor NOR2_1929 (G5114gat, G5059gat, G4995gat);
nor NOR2_1930 (G5115gat, G5063gat, G5064gat);
nor NOR2_1931 (G5118gat, G5065gat, G5066gat);
nor NOR2_1932 (G5121gat, G5067gat, G5068gat);
nor NOR2_1933 (G5124gat, G5069gat, G5070gat);
nor NOR2_1934 (G5127gat, G5071gat, G5072gat);
nor NOR2_1935 (G5130gat, G5073gat, G771gat);
nor NOR2_1936 (G5134gat, G5023gat, G5076gat);
nor NOR2_1937 (G5135gat, G5076gat, G819gat);
nor NOR2_1938 (G5136gat, G4907gat, G5076gat);
nor NOR2_1939 (G5139gat, G5080gat, G5081gat);
nor NOR2_1940 (G5142gat, G5085gat, G5082gat);
nor NOR2_1941 (G5146gat, G5035gat, G5088gat);
nor NOR2_1942 (G5147gat, G5088gat, G5032gat);
nor NOR2_1943 (G5148gat, G5092gat, G5093gat);
nor NOR2_1944 (G5151gat, G5094gat, G1014gat);
nor NOR2_1945 (G5155gat, G5044gat, G5097gat);
nor NOR2_1946 (G5156gat, G5097gat, G1062gat);
nor NOR2_1947 (G5157gat, G4928gat, G5097gat);
nor NOR2_1948 (G5160gat, G5101gat, G5102gat);
nor NOR2_1949 (G5163gat, G5106gat, G5103gat);
nor NOR2_1950 (G5167gat, G5056gat, G5109gat);
nor NOR2_1951 (G5168gat, G5109gat, G5053gat);
nor NOR2_1952 (G5169gat, G5113gat, G5114gat);
nor NOR2_1953 (G5172gat, G5115gat, G1257gat);
nor NOR2_1954 (G5176gat, G5118gat, G579gat);
nor NOR2_1955 (G5180gat, G5121gat, G627gat);
nor NOR2_1956 (G5184gat, G5124gat, G675gat);
nor NOR2_1957 (G5188gat, G5127gat, G723gat);
nor NOR2_1958 (G5192gat, G5073gat, G5130gat);
nor NOR2_1959 (G5193gat, G5130gat, G771gat);
nor NOR2_1960 (G5194gat, G4959gat, G5130gat);
nor NOR2_1961 (G5197gat, G5134gat, G5135gat);
nor NOR2_1962 (G5200gat, G5139gat, G5136gat);
nor NOR2_1963 (G5204gat, G5085gat, G5142gat);
nor NOR2_1964 (G5205gat, G5142gat, G5082gat);
nor NOR2_1965 (G5206gat, G5146gat, G5147gat);
nor NOR2_1966 (G5209gat, G5148gat, G966gat);
nor NOR2_1967 (G5213gat, G5094gat, G5151gat);
nor NOR2_1968 (G5214gat, G5151gat, G1014gat);
nor NOR2_1969 (G5215gat, G4980gat, G5151gat);
nor NOR2_1970 (G5218gat, G5155gat, G5156gat);
nor NOR2_1971 (G5221gat, G5160gat, G5157gat);
nor NOR2_1972 (G5225gat, G5106gat, G5163gat);
nor NOR2_1973 (G5226gat, G5163gat, G5103gat);
nor NOR2_1974 (G5227gat, G5167gat, G5168gat);
nor NOR2_1975 (G5230gat, G5169gat, G1209gat);
nor NOR2_1976 (G5234gat, G5115gat, G5172gat);
nor NOR2_1977 (G5235gat, G5172gat, G1257gat);
nor NOR2_1978 (G5236gat, G5001gat, G5172gat);
nor NOR2_1979 (G5239gat, G5118gat, G5176gat);
nor NOR2_1980 (G5240gat, G5176gat, G579gat);
nor NOR2_1981 (G5241gat, G5005gat, G5176gat);
nor NOR2_1982 (G5244gat, G5121gat, G5180gat);
nor NOR2_1983 (G5245gat, G5180gat, G627gat);
nor NOR2_1984 (G5246gat, G5009gat, G5180gat);
nor NOR2_1985 (G5249gat, G5124gat, G5184gat);
nor NOR2_1986 (G5250gat, G5184gat, G675gat);
nor NOR2_1987 (G5251gat, G5013gat, G5184gat);
nor NOR2_1988 (G5254gat, G5127gat, G5188gat);
nor NOR2_1989 (G5255gat, G5188gat, G723gat);
nor NOR2_1990 (G5256gat, G5017gat, G5188gat);
nor NOR2_1991 (G5259gat, G5192gat, G5193gat);
nor NOR2_1992 (G5262gat, G5197gat, G5194gat);
nor NOR2_1993 (G5266gat, G5139gat, G5200gat);
nor NOR2_1994 (G5267gat, G5200gat, G5136gat);
nor NOR2_1995 (G5268gat, G5204gat, G5205gat);
nor NOR2_1996 (G5271gat, G5206gat, G918gat);
nor NOR2_1997 (G5275gat, G5148gat, G5209gat);
nor NOR2_1998 (G5276gat, G5209gat, G966gat);
nor NOR2_1999 (G5277gat, G5038gat, G5209gat);
nor NOR2_2000 (G5280gat, G5213gat, G5214gat);
nor NOR2_2001 (G5283gat, G5218gat, G5215gat);
nor NOR2_2002 (G5287gat, G5160gat, G5221gat);
nor NOR2_2003 (G5288gat, G5221gat, G5157gat);
nor NOR2_2004 (G5289gat, G5225gat, G5226gat);
nor NOR2_2005 (G5292gat, G5227gat, G1161gat);
nor NOR2_2006 (G5296gat, G5169gat, G5230gat);
nor NOR2_2007 (G5297gat, G5230gat, G1209gat);
nor NOR2_2008 (G5298gat, G5059gat, G5230gat);
nor NOR2_2009 (G5301gat, G5234gat, G5235gat);
nor NOR2_2010 (G5304gat, G1305gat, G5236gat);
nor NOR2_2011 (G5308gat, G5239gat, G5240gat);
nor NOR2_2012 (G5309gat, G5244gat, G5245gat);
nor NOR2_2013 (G5312gat, G5249gat, G5250gat);
nor NOR2_2014 (G5315gat, G5254gat, G5255gat);
nor NOR2_2015 (G5318gat, G5259gat, G5256gat);
nor NOR2_2016 (G5322gat, G5197gat, G5262gat);
nor NOR2_2017 (G5323gat, G5262gat, G5194gat);
nor NOR2_2018 (G5324gat, G5266gat, G5267gat);
nor NOR2_2019 (G5327gat, G5268gat, G870gat);
nor NOR2_2020 (G5331gat, G5206gat, G5271gat);
nor NOR2_2021 (G5332gat, G5271gat, G918gat);
nor NOR2_2022 (G5333gat, G5088gat, G5271gat);
nor NOR2_2023 (G5336gat, G5275gat, G5276gat);
nor NOR2_2024 (G5339gat, G5280gat, G5277gat);
nor NOR2_2025 (G5343gat, G5218gat, G5283gat);
nor NOR2_2026 (G5344gat, G5283gat, G5215gat);
nor NOR2_2027 (G5345gat, G5287gat, G5288gat);
nor NOR2_2028 (G5348gat, G5289gat, G1113gat);
nor NOR2_2029 (G5352gat, G5227gat, G5292gat);
nor NOR2_2030 (G5353gat, G5292gat, G1161gat);
nor NOR2_2031 (G5354gat, G5109gat, G5292gat);
nor NOR2_2032 (G5357gat, G5296gat, G5297gat);
nor NOR2_2033 (G5360gat, G5301gat, G5298gat);
nor NOR2_2034 (G5364gat, G1305gat, G5304gat);
nor NOR2_2035 (G5365gat, G5304gat, G5236gat);
nor NOR2_2036 (G5366gat, G5309gat, G5241gat);
nor NOR2_2037 (G5370gat, G5312gat, G5246gat);
nor NOR2_2038 (G5374gat, G5315gat, G5251gat);
nor NOR2_2039 (G5378gat, G5259gat, G5318gat);
nor NOR2_2040 (G5379gat, G5318gat, G5256gat);
nor NOR2_2041 (G5380gat, G5322gat, G5323gat);
nor NOR2_2042 (G5383gat, G5324gat, G822gat);
nor NOR2_2043 (G5387gat, G5268gat, G5327gat);
nor NOR2_2044 (G5388gat, G5327gat, G870gat);
nor NOR2_2045 (G5389gat, G5142gat, G5327gat);
nor NOR2_2046 (G5392gat, G5331gat, G5332gat);
nor NOR2_2047 (G5395gat, G5336gat, G5333gat);
nor NOR2_2048 (G5399gat, G5280gat, G5339gat);
nor NOR2_2049 (G5400gat, G5339gat, G5277gat);
nor NOR2_2050 (G5401gat, G5343gat, G5344gat);
nor NOR2_2051 (G5404gat, G5345gat, G1065gat);
nor NOR2_2052 (G5408gat, G5289gat, G5348gat);
nor NOR2_2053 (G5409gat, G5348gat, G1113gat);
nor NOR2_2054 (G5410gat, G5163gat, G5348gat);
nor NOR2_2055 (G5413gat, G5352gat, G5353gat);
nor NOR2_2056 (G5416gat, G5357gat, G5354gat);
nor NOR2_2057 (G5420gat, G5301gat, G5360gat);
nor NOR2_2058 (G5421gat, G5360gat, G5298gat);
nor NOR2_2059 (G5422gat, G5364gat, G5365gat);
nor NOR2_2060 (G5425gat, G5309gat, G5366gat);
nor NOR2_2061 (G5426gat, G5366gat, G5241gat);
nor NOR2_2062 (G5427gat, G5312gat, G5370gat);
nor NOR2_2063 (G5428gat, G5370gat, G5246gat);
nor NOR2_2064 (G5429gat, G5315gat, G5374gat);
nor NOR2_2065 (G5430gat, G5374gat, G5251gat);
nor NOR2_2066 (G5431gat, G5378gat, G5379gat);
nor NOR2_2067 (G5434gat, G5380gat, G774gat);
nor NOR2_2068 (G5438gat, G5324gat, G5383gat);
nor NOR2_2069 (G5439gat, G5383gat, G822gat);
nor NOR2_2070 (G5440gat, G5200gat, G5383gat);
nor NOR2_2071 (G5443gat, G5387gat, G5388gat);
nor NOR2_2072 (G5446gat, G5392gat, G5389gat);
nor NOR2_2073 (G5450gat, G5336gat, G5395gat);
nor NOR2_2074 (G5451gat, G5395gat, G5333gat);
nor NOR2_2075 (G5452gat, G5399gat, G5400gat);
nor NOR2_2076 (G5455gat, G5401gat, G1017gat);
nor NOR2_2077 (G5459gat, G5345gat, G5404gat);
nor NOR2_2078 (G5460gat, G5404gat, G1065gat);
nor NOR2_2079 (G5461gat, G5221gat, G5404gat);
nor NOR2_2080 (G5464gat, G5408gat, G5409gat);
nor NOR2_2081 (G5467gat, G5413gat, G5410gat);
nor NOR2_2082 (G5471gat, G5357gat, G5416gat);
nor NOR2_2083 (G5472gat, G5416gat, G5354gat);
nor NOR2_2084 (G5473gat, G5420gat, G5421gat);
nor NOR2_2085 (G5476gat, G5422gat, G1260gat);
nor NOR2_2086 (G5480gat, G5425gat, G5426gat);
nor NOR2_2087 (G5483gat, G5427gat, G5428gat);
nor NOR2_2088 (G5486gat, G5429gat, G5430gat);
nor NOR2_2089 (G5489gat, G5431gat, G726gat);
nor NOR2_2090 (G5493gat, G5380gat, G5434gat);
nor NOR2_2091 (G5494gat, G5434gat, G774gat);
nor NOR2_2092 (G5495gat, G5262gat, G5434gat);
nor NOR2_2093 (G5498gat, G5438gat, G5439gat);
nor NOR2_2094 (G5501gat, G5443gat, G5440gat);
nor NOR2_2095 (G5505gat, G5392gat, G5446gat);
nor NOR2_2096 (G5506gat, G5446gat, G5389gat);
nor NOR2_2097 (G5507gat, G5450gat, G5451gat);
nor NOR2_2098 (G5510gat, G5452gat, G969gat);
nor NOR2_2099 (G5514gat, G5401gat, G5455gat);
nor NOR2_2100 (G5515gat, G5455gat, G1017gat);
nor NOR2_2101 (G5516gat, G5283gat, G5455gat);
nor NOR2_2102 (G5519gat, G5459gat, G5460gat);
nor NOR2_2103 (G5522gat, G5464gat, G5461gat);
nor NOR2_2104 (G5526gat, G5413gat, G5467gat);
nor NOR2_2105 (G5527gat, G5467gat, G5410gat);
nor NOR2_2106 (G5528gat, G5471gat, G5472gat);
nor NOR2_2107 (G5531gat, G5473gat, G1212gat);
nor NOR2_2108 (G5535gat, G5422gat, G5476gat);
nor NOR2_2109 (G5536gat, G5476gat, G1260gat);
nor NOR2_2110 (G5537gat, G5304gat, G5476gat);
nor NOR2_2111 (G5540gat, G5480gat, G582gat);
nor NOR2_2112 (G5544gat, G5483gat, G630gat);
nor NOR2_2113 (G5548gat, G5486gat, G678gat);
nor NOR2_2114 (G5552gat, G5431gat, G5489gat);
nor NOR2_2115 (G5553gat, G5489gat, G726gat);
nor NOR2_2116 (G5554gat, G5318gat, G5489gat);
nor NOR2_2117 (G5557gat, G5493gat, G5494gat);
nor NOR2_2118 (G5560gat, G5498gat, G5495gat);
nor NOR2_2119 (G5564gat, G5443gat, G5501gat);
nor NOR2_2120 (G5565gat, G5501gat, G5440gat);
nor NOR2_2121 (G5566gat, G5505gat, G5506gat);
nor NOR2_2122 (G5569gat, G5507gat, G921gat);
nor NOR2_2123 (G5573gat, G5452gat, G5510gat);
nor NOR2_2124 (G5574gat, G5510gat, G969gat);
nor NOR2_2125 (G5575gat, G5339gat, G5510gat);
nor NOR2_2126 (G5578gat, G5514gat, G5515gat);
nor NOR2_2127 (G5581gat, G5519gat, G5516gat);
nor NOR2_2128 (G5585gat, G5464gat, G5522gat);
nor NOR2_2129 (G5586gat, G5522gat, G5461gat);
nor NOR2_2130 (G5587gat, G5526gat, G5527gat);
nor NOR2_2131 (G5590gat, G5528gat, G1164gat);
nor NOR2_2132 (G5594gat, G5473gat, G5531gat);
nor NOR2_2133 (G5595gat, G5531gat, G1212gat);
nor NOR2_2134 (G5596gat, G5360gat, G5531gat);
nor NOR2_2135 (G5599gat, G5535gat, G5536gat);
nor NOR2_2136 (G5602gat, G1308gat, G5537gat);
nor NOR2_2137 (G5606gat, G5480gat, G5540gat);
nor NOR2_2138 (G5607gat, G5540gat, G582gat);
nor NOR2_2139 (G5608gat, G5366gat, G5540gat);
nor NOR2_2140 (G5611gat, G5483gat, G5544gat);
nor NOR2_2141 (G5612gat, G5544gat, G630gat);
nor NOR2_2142 (G5613gat, G5370gat, G5544gat);
nor NOR2_2143 (G5616gat, G5486gat, G5548gat);
nor NOR2_2144 (G5617gat, G5548gat, G678gat);
nor NOR2_2145 (G5618gat, G5374gat, G5548gat);
nor NOR2_2146 (G5621gat, G5552gat, G5553gat);
nor NOR2_2147 (G5624gat, G5557gat, G5554gat);
nor NOR2_2148 (G5628gat, G5498gat, G5560gat);
nor NOR2_2149 (G5629gat, G5560gat, G5495gat);
nor NOR2_2150 (G5630gat, G5564gat, G5565gat);
nor NOR2_2151 (G5633gat, G5566gat, G873gat);
nor NOR2_2152 (G5637gat, G5507gat, G5569gat);
nor NOR2_2153 (G5638gat, G5569gat, G921gat);
nor NOR2_2154 (G5639gat, G5395gat, G5569gat);
nor NOR2_2155 (G5642gat, G5573gat, G5574gat);
nor NOR2_2156 (G5645gat, G5578gat, G5575gat);
nor NOR2_2157 (G5649gat, G5519gat, G5581gat);
nor NOR2_2158 (G5650gat, G5581gat, G5516gat);
nor NOR2_2159 (G5651gat, G5585gat, G5586gat);
nor NOR2_2160 (G5654gat, G5587gat, G1116gat);
nor NOR2_2161 (G5658gat, G5528gat, G5590gat);
nor NOR2_2162 (G5659gat, G5590gat, G1164gat);
nor NOR2_2163 (G5660gat, G5416gat, G5590gat);
nor NOR2_2164 (G5663gat, G5594gat, G5595gat);
nor NOR2_2165 (G5666gat, G5599gat, G5596gat);
nor NOR2_2166 (G5670gat, G1308gat, G5602gat);
nor NOR2_2167 (G5671gat, G5602gat, G5537gat);
nor NOR2_2168 (G5672gat, G5606gat, G5607gat);
nor NOR2_2169 (G5673gat, G5611gat, G5612gat);
nor NOR2_2170 (G5676gat, G5616gat, G5617gat);
nor NOR2_2171 (G5679gat, G5621gat, G5618gat);
nor NOR2_2172 (G5683gat, G5557gat, G5624gat);
nor NOR2_2173 (G5684gat, G5624gat, G5554gat);
nor NOR2_2174 (G5685gat, G5628gat, G5629gat);
nor NOR2_2175 (G5688gat, G5630gat, G825gat);
nor NOR2_2176 (G5692gat, G5566gat, G5633gat);
nor NOR2_2177 (G5693gat, G5633gat, G873gat);
nor NOR2_2178 (G5694gat, G5446gat, G5633gat);
nor NOR2_2179 (G5697gat, G5637gat, G5638gat);
nor NOR2_2180 (G5700gat, G5642gat, G5639gat);
nor NOR2_2181 (G5704gat, G5578gat, G5645gat);
nor NOR2_2182 (G5705gat, G5645gat, G5575gat);
nor NOR2_2183 (G5706gat, G5649gat, G5650gat);
nor NOR2_2184 (G5709gat, G5651gat, G1068gat);
nor NOR2_2185 (G5713gat, G5587gat, G5654gat);
nor NOR2_2186 (G5714gat, G5654gat, G1116gat);
nor NOR2_2187 (G5715gat, G5467gat, G5654gat);
nor NOR2_2188 (G5718gat, G5658gat, G5659gat);
nor NOR2_2189 (G5721gat, G5663gat, G5660gat);
nor NOR2_2190 (G5725gat, G5599gat, G5666gat);
nor NOR2_2191 (G5726gat, G5666gat, G5596gat);
nor NOR2_2192 (G5727gat, G5670gat, G5671gat);
nor NOR2_2193 (G5730gat, G5673gat, G5608gat);
nor NOR2_2194 (G5734gat, G5676gat, G5613gat);
nor NOR2_2195 (G5738gat, G5621gat, G5679gat);
nor NOR2_2196 (G5739gat, G5679gat, G5618gat);
nor NOR2_2197 (G5740gat, G5683gat, G5684gat);
nor NOR2_2198 (G5743gat, G5685gat, G777gat);
nor NOR2_2199 (G5747gat, G5630gat, G5688gat);
nor NOR2_2200 (G5748gat, G5688gat, G825gat);
nor NOR2_2201 (G5749gat, G5501gat, G5688gat);
nor NOR2_2202 (G5752gat, G5692gat, G5693gat);
nor NOR2_2203 (G5755gat, G5697gat, G5694gat);
nor NOR2_2204 (G5759gat, G5642gat, G5700gat);
nor NOR2_2205 (G5760gat, G5700gat, G5639gat);
nor NOR2_2206 (G5761gat, G5704gat, G5705gat);
nor NOR2_2207 (G5764gat, G5706gat, G1020gat);
nor NOR2_2208 (G5768gat, G5651gat, G5709gat);
nor NOR2_2209 (G5769gat, G5709gat, G1068gat);
nor NOR2_2210 (G5770gat, G5522gat, G5709gat);
nor NOR2_2211 (G5773gat, G5713gat, G5714gat);
nor NOR2_2212 (G5776gat, G5718gat, G5715gat);
nor NOR2_2213 (G5780gat, G5663gat, G5721gat);
nor NOR2_2214 (G5781gat, G5721gat, G5660gat);
nor NOR2_2215 (G5782gat, G5725gat, G5726gat);
nor NOR2_2216 (G5785gat, G5673gat, G5730gat);
nor NOR2_2217 (G5786gat, G5730gat, G5608gat);
nor NOR2_2218 (G5787gat, G5676gat, G5734gat);
nor NOR2_2219 (G5788gat, G5734gat, G5613gat);
nor NOR2_2220 (G5789gat, G5738gat, G5739gat);
nor NOR2_2221 (G5792gat, G5740gat, G729gat);
nor NOR2_2222 (G5796gat, G5685gat, G5743gat);
nor NOR2_2223 (G5797gat, G5743gat, G777gat);
nor NOR2_2224 (G5798gat, G5560gat, G5743gat);
nor NOR2_2225 (G5801gat, G5747gat, G5748gat);
nor NOR2_2226 (G5804gat, G5752gat, G5749gat);
nor NOR2_2227 (G5808gat, G5697gat, G5755gat);
nor NOR2_2228 (G5809gat, G5755gat, G5694gat);
nor NOR2_2229 (G5810gat, G5759gat, G5760gat);
nor NOR2_2230 (G5813gat, G5761gat, G972gat);
nor NOR2_2231 (G5817gat, G5706gat, G5764gat);
nor NOR2_2232 (G5818gat, G5764gat, G1020gat);
nor NOR2_2233 (G5819gat, G5581gat, G5764gat);
nor NOR2_2234 (G5822gat, G5768gat, G5769gat);
nor NOR2_2235 (G5825gat, G5773gat, G5770gat);
nor NOR2_2236 (G5829gat, G5718gat, G5776gat);
nor NOR2_2237 (G5830gat, G5776gat, G5715gat);
nor NOR2_2238 (G5831gat, G5780gat, G5781gat);
nor NOR2_2239 (G5834gat, G5785gat, G5786gat);
nor NOR2_2240 (G5837gat, G5787gat, G5788gat);
nor NOR2_2241 (G5840gat, G5789gat, G681gat);
nor NOR2_2242 (G5844gat, G5740gat, G5792gat);
nor NOR2_2243 (G5845gat, G5792gat, G729gat);
nor NOR2_2244 (G5846gat, G5624gat, G5792gat);
nor NOR2_2245 (G5849gat, G5796gat, G5797gat);
nor NOR2_2246 (G5852gat, G5801gat, G5798gat);
nor NOR2_2247 (G5856gat, G5752gat, G5804gat);
nor NOR2_2248 (G5857gat, G5804gat, G5749gat);
nor NOR2_2249 (G5858gat, G5808gat, G5809gat);
nor NOR2_2250 (G5861gat, G5810gat, G924gat);
nor NOR2_2251 (G5865gat, G5761gat, G5813gat);
nor NOR2_2252 (G5866gat, G5813gat, G972gat);
nor NOR2_2253 (G5867gat, G5645gat, G5813gat);
nor NOR2_2254 (G5870gat, G5817gat, G5818gat);
nor NOR2_2255 (G5873gat, G5822gat, G5819gat);
nor NOR2_2256 (G5877gat, G5773gat, G5825gat);
nor NOR2_2257 (G5878gat, G5825gat, G5770gat);
nor NOR2_2258 (G5879gat, G5829gat, G5830gat);
nor NOR2_2259 (G5882gat, G5834gat, G585gat);
nor NOR2_2260 (G5886gat, G5837gat, G633gat);
nor NOR2_2261 (G5890gat, G5789gat, G5840gat);
nor NOR2_2262 (G5891gat, G5840gat, G681gat);
nor NOR2_2263 (G5892gat, G5679gat, G5840gat);
nor NOR2_2264 (G5895gat, G5844gat, G5845gat);
nor NOR2_2265 (G5898gat, G5849gat, G5846gat);
nor NOR2_2266 (G5902gat, G5801gat, G5852gat);
nor NOR2_2267 (G5903gat, G5852gat, G5798gat);
nor NOR2_2268 (G5904gat, G5856gat, G5857gat);
nor NOR2_2269 (G5907gat, G5858gat, G876gat);
nor NOR2_2270 (G5911gat, G5810gat, G5861gat);
nor NOR2_2271 (G5912gat, G5861gat, G924gat);
nor NOR2_2272 (G5913gat, G5700gat, G5861gat);
nor NOR2_2273 (G5916gat, G5865gat, G5866gat);
nor NOR2_2274 (G5919gat, G5870gat, G5867gat);
nor NOR2_2275 (G5923gat, G5822gat, G5873gat);
nor NOR2_2276 (G5924gat, G5873gat, G5819gat);
nor NOR2_2277 (G5925gat, G5877gat, G5878gat);
nor NOR2_2278 (G5928gat, G5834gat, G5882gat);
nor NOR2_2279 (G5929gat, G5882gat, G585gat);
nor NOR2_2280 (G5930gat, G5730gat, G5882gat);
nor NOR2_2281 (G5933gat, G5837gat, G5886gat);
nor NOR2_2282 (G5934gat, G5886gat, G633gat);
nor NOR2_2283 (G5935gat, G5734gat, G5886gat);
nor NOR2_2284 (G5938gat, G5890gat, G5891gat);
nor NOR2_2285 (G5941gat, G5895gat, G5892gat);
nor NOR2_2286 (G5945gat, G5849gat, G5898gat);
nor NOR2_2287 (G5946gat, G5898gat, G5846gat);
nor NOR2_2288 (G5947gat, G5902gat, G5903gat);
nor NOR2_2289 (G5950gat, G5904gat, G828gat);
nor NOR2_2290 (G5954gat, G5858gat, G5907gat);
nor NOR2_2291 (G5955gat, G5907gat, G876gat);
nor NOR2_2292 (G5956gat, G5755gat, G5907gat);
nor NOR2_2293 (G5959gat, G5911gat, G5912gat);
nor NOR2_2294 (G5962gat, G5916gat, G5913gat);
nor NOR2_2295 (G5966gat, G5870gat, G5919gat);
nor NOR2_2296 (G5967gat, G5919gat, G5867gat);
nor NOR2_2297 (G5968gat, G5923gat, G5924gat);
nor NOR2_2298 (G5971gat, G5928gat, G5929gat);
nor NOR2_2299 (G5972gat, G5933gat, G5934gat);
nor NOR2_2300 (G5975gat, G5938gat, G5935gat);
nor NOR2_2301 (G5979gat, G5895gat, G5941gat);
nor NOR2_2302 (G5980gat, G5941gat, G5892gat);
nor NOR2_2303 (G5981gat, G5945gat, G5946gat);
nor NOR2_2304 (G5984gat, G5947gat, G780gat);
nor NOR2_2305 (G5988gat, G5904gat, G5950gat);
nor NOR2_2306 (G5989gat, G5950gat, G828gat);
nor NOR2_2307 (G5990gat, G5804gat, G5950gat);
nor NOR2_2308 (G5993gat, G5954gat, G5955gat);
nor NOR2_2309 (G5996gat, G5959gat, G5956gat);
nor NOR2_2310 (G6000gat, G5916gat, G5962gat);
nor NOR2_2311 (G6001gat, G5962gat, G5913gat);
nor NOR2_2312 (G6002gat, G5966gat, G5967gat);
nor NOR2_2313 (G6005gat, G5972gat, G5930gat);
nor NOR2_2314 (G6009gat, G5938gat, G5975gat);
nor NOR2_2315 (G6010gat, G5975gat, G5935gat);
nor NOR2_2316 (G6011gat, G5979gat, G5980gat);
nor NOR2_2317 (G6014gat, G5981gat, G732gat);
nor NOR2_2318 (G6018gat, G5947gat, G5984gat);
nor NOR2_2319 (G6019gat, G5984gat, G780gat);
nor NOR2_2320 (G6020gat, G5852gat, G5984gat);
nor NOR2_2321 (G6023gat, G5988gat, G5989gat);
nor NOR2_2322 (G6026gat, G5993gat, G5990gat);
nor NOR2_2323 (G6030gat, G5959gat, G5996gat);
nor NOR2_2324 (G6031gat, G5996gat, G5956gat);
nor NOR2_2325 (G6032gat, G6000gat, G6001gat);
nor NOR2_2326 (G6035gat, G5972gat, G6005gat);
nor NOR2_2327 (G6036gat, G6005gat, G5930gat);
nor NOR2_2328 (G6037gat, G6009gat, G6010gat);
nor NOR2_2329 (G6040gat, G6011gat, G684gat);
nor NOR2_2330 (G6044gat, G5981gat, G6014gat);
nor NOR2_2331 (G6045gat, G6014gat, G732gat);
nor NOR2_2332 (G6046gat, G5898gat, G6014gat);
nor NOR2_2333 (G6049gat, G6018gat, G6019gat);
nor NOR2_2334 (G6052gat, G6023gat, G6020gat);
nor NOR2_2335 (G6056gat, G5993gat, G6026gat);
nor NOR2_2336 (G6057gat, G6026gat, G5990gat);
nor NOR2_2337 (G6058gat, G6030gat, G6031gat);
nor NOR2_2338 (G6061gat, G6035gat, G6036gat);
nor NOR2_2339 (G6064gat, G6037gat, G636gat);
nor NOR2_2340 (G6068gat, G6011gat, G6040gat);
nor NOR2_2341 (G6069gat, G6040gat, G684gat);
nor NOR2_2342 (G6070gat, G5941gat, G6040gat);
nor NOR2_2343 (G6073gat, G6044gat, G6045gat);
nor NOR2_2344 (G6076gat, G6049gat, G6046gat);
nor NOR2_2345 (G6080gat, G6023gat, G6052gat);
nor NOR2_2346 (G6081gat, G6052gat, G6020gat);
nor NOR2_2347 (G6082gat, G6056gat, G6057gat);
nor NOR2_2348 (G6085gat, G6061gat, G588gat);
nor NOR2_2349 (G6089gat, G6037gat, G6064gat);
nor NOR2_2350 (G6090gat, G6064gat, G636gat);
nor NOR2_2351 (G6091gat, G5975gat, G6064gat);
nor NOR2_2352 (G6094gat, G6068gat, G6069gat);
nor NOR2_2353 (G6097gat, G6073gat, G6070gat);
nor NOR2_2354 (G6101gat, G6049gat, G6076gat);
nor NOR2_2355 (G6102gat, G6076gat, G6046gat);
nor NOR2_2356 (G6103gat, G6080gat, G6081gat);
nor NOR2_2357 (G6106gat, G6061gat, G6085gat);
nor NOR2_2358 (G6107gat, G6085gat, G588gat);
nor NOR2_2359 (G6108gat, G6005gat, G6085gat);
nor NOR2_2360 (G6111gat, G6089gat, G6090gat);
nor NOR2_2361 (G6114gat, G6094gat, G6091gat);
nor NOR2_2362 (G6118gat, G6073gat, G6097gat);
nor NOR2_2363 (G6119gat, G6097gat, G6070gat);
nor NOR2_2364 (G6120gat, G6101gat, G6102gat);
nor NOR2_2365 (G6123gat, G6106gat, G6107gat);
nor NOR2_2366 (G6124gat, G6111gat, G6108gat);
nor NOR2_2367 (G6128gat, G6094gat, G6114gat);
nor NOR2_2368 (G6129gat, G6114gat, G6091gat);
nor NOR2_2369 (G6130gat, G6118gat, G6119gat);
nor NOR2_2370 (G6133gat, G6111gat, G6124gat);
nor NOR2_2371 (G6134gat, G6124gat, G6108gat);
nor NOR2_2372 (G6135gat, G6128gat, G6129gat);
nor NOR2_2373 (G6138gat, G6133gat, G6134gat);
not NOT1_2374 (G6141gat, G6138gat);
nor NOR2_2375 (G6145gat, G6138gat, G6141gat);
not NOT1_2376 (G6146gat, G6141gat);
nor NOR2_2377 (G6147gat, G6124gat, G6141gat);
nor NOR2_2378 (G6150gat, G6145gat, G6146gat);
nor NOR2_2379 (G6151gat, G6135gat, G6147gat);
nor NOR2_2380 (G6155gat, G6135gat, G6151gat);
nor NOR2_2381 (G6156gat, G6151gat, G6147gat);
nor NOR2_2382 (G6157gat, G6114gat, G6151gat);
nor NOR2_2383 (G6160gat, G6155gat, G6156gat);
nor NOR2_2384 (G6161gat, G6130gat, G6157gat);
nor NOR2_2385 (G6165gat, G6130gat, G6161gat);
nor NOR2_2386 (G6166gat, G6161gat, G6157gat);
nor NOR2_2387 (G6167gat, G6097gat, G6161gat);
nor NOR2_2388 (G6170gat, G6165gat, G6166gat);
nor NOR2_2389 (G6171gat, G6120gat, G6167gat);
nor NOR2_2390 (G6175gat, G6120gat, G6171gat);
nor NOR2_2391 (G6176gat, G6171gat, G6167gat);
nor NOR2_2392 (G6177gat, G6076gat, G6171gat);
nor NOR2_2393 (G6180gat, G6175gat, G6176gat);
nor NOR2_2394 (G6181gat, G6103gat, G6177gat);
nor NOR2_2395 (G6185gat, G6103gat, G6181gat);
nor NOR2_2396 (G6186gat, G6181gat, G6177gat);
nor NOR2_2397 (G6187gat, G6052gat, G6181gat);
nor NOR2_2398 (G6190gat, G6185gat, G6186gat);
nor NOR2_2399 (G6191gat, G6082gat, G6187gat);
nor NOR2_2400 (G6195gat, G6082gat, G6191gat);
nor NOR2_2401 (G6196gat, G6191gat, G6187gat);
nor NOR2_2402 (G6197gat, G6026gat, G6191gat);
nor NOR2_2403 (G6200gat, G6195gat, G6196gat);
nor NOR2_2404 (G6201gat, G6058gat, G6197gat);
nor NOR2_2405 (G6205gat, G6058gat, G6201gat);
nor NOR2_2406 (G6206gat, G6201gat, G6197gat);
nor NOR2_2407 (G6207gat, G5996gat, G6201gat);
nor NOR2_2408 (G6210gat, G6205gat, G6206gat);
nor NOR2_2409 (G6211gat, G6032gat, G6207gat);
nor NOR2_2410 (G6215gat, G6032gat, G6211gat);
nor NOR2_2411 (G6216gat, G6211gat, G6207gat);
nor NOR2_2412 (G6217gat, G5962gat, G6211gat);
nor NOR2_2413 (G6220gat, G6215gat, G6216gat);
nor NOR2_2414 (G6221gat, G6002gat, G6217gat);
nor NOR2_2415 (G6225gat, G6002gat, G6221gat);
nor NOR2_2416 (G6226gat, G6221gat, G6217gat);
nor NOR2_2417 (G6227gat, G5919gat, G6221gat);
nor NOR2_2418 (G6230gat, G6225gat, G6226gat);
nor NOR2_2419 (G6231gat, G5968gat, G6227gat);
nor NOR2_2420 (G6235gat, G5968gat, G6231gat);
nor NOR2_2421 (G6236gat, G6231gat, G6227gat);
nor NOR2_2422 (G6237gat, G5873gat, G6231gat);
nor NOR2_2423 (G6240gat, G6235gat, G6236gat);
nor NOR2_2424 (G6241gat, G5925gat, G6237gat);
nor NOR2_2425 (G6245gat, G5925gat, G6241gat);
nor NOR2_2426 (G6246gat, G6241gat, G6237gat);
nor NOR2_2427 (G6247gat, G5825gat, G6241gat);
nor NOR2_2428 (G6250gat, G6245gat, G6246gat);
nor NOR2_2429 (G6251gat, G5879gat, G6247gat);
nor NOR2_2430 (G6255gat, G5879gat, G6251gat);
nor NOR2_2431 (G6256gat, G6251gat, G6247gat);
nor NOR2_2432 (G6257gat, G5776gat, G6251gat);
nor NOR2_2433 (G6260gat, G6255gat, G6256gat);
nor NOR2_2434 (G6261gat, G5831gat, G6257gat);
nor NOR2_2435 (G6265gat, G5831gat, G6261gat);
nor NOR2_2436 (G6266gat, G6261gat, G6257gat);
nor NOR2_2437 (G6267gat, G5721gat, G6261gat);
nor NOR2_2438 (G6270gat, G6265gat, G6266gat);
nor NOR2_2439 (G6271gat, G5782gat, G6267gat);
nor NOR2_2440 (G6275gat, G5782gat, G6271gat);
nor NOR2_2441 (G6276gat, G6271gat, G6267gat);
nor NOR2_2442 (G6277gat, G5666gat, G6271gat);
nor NOR2_2443 (G6280gat, G6275gat, G6276gat);
nor NOR2_2444 (G6281gat, G5727gat, G6277gat);
nor NOR2_2445 (G6285gat, G5727gat, G6281gat);
nor NOR2_2446 (G6286gat, G6281gat, G6277gat);
nor NOR2_2447 (G6287gat, G5602gat, G6281gat);
nor NOR2_2448 (G6288gat, G6285gat, G6286gat);

endmodule