module DFF(Q, clk, D);
input D;
input clk;
output Q;
always @(clk)
begin
  Q <= D;
end
endmodule


module c1355_libar_8k(G1gat,G8gat,G15gat,G22gat,G29gat,G36gat,G43gat,G50gat,G57gat,G64gat,G71gat,G78gat,G85gat,G92gat,G99gat,G106gat,G113gat,G120gat,G127gat,G134gat,G141gat,G148gat,G155gat,G162gat,G169gat,G176gat,G183gat,G190gat,G197gat,G204gat,G211gat,G218gat,G225gat,G226gat,G227gat,G228gat,G229gat,G230gat,G231gat,G232gat,G233gat,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,G1324gat,G1325gat,G1326gat,G1327gat,G1328gat,G1329gat,G1330gat,G1331gat,G1332gat,G1333gat,G1334gat,G1335gat,G1336gat,G1337gat,G1338gat,G1339gat,G1340gat,G1341gat,G1342gat,G1343gat,G1344gat,G1345gat,G1346gat,G1347gat,G1348gat,G1349gat,G1350gat,G1351gat,G1352gat,G1353gat,G1354gat,G1355gat);

input G1gat,G8gat,G15gat,G22gat,G29gat,G36gat,G43gat,G50gat,G57gat,G64gat,G71gat,G78gat,G85gat,G92gat,G99gat,G106gat,G113gat,G120gat,G127gat,G134gat,G141gat,G148gat,G155gat,G162gat,G169gat,G176gat,G183gat,G190gat,G197gat,G204gat,G211gat,G218gat,G225gat,G226gat,G227gat,G228gat,G229gat,G230gat,G231gat,G232gat,G233gat,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7;
output G1324gat,G1325gat,G1326gat,G1327gat,G1328gat,G1329gat,G1330gat,G1331gat,G1332gat,G1333gat,G1334gat,G1335gat,G1336gat,G1337gat,G1338gat,G1339gat,G1340gat,G1341gat,G1342gat,G1343gat,G1344gat,G1345gat,G1346gat,G1347gat,G1348gat,G1349gat,G1350gat,G1351gat,G1352gat,G1353gat,G1354gat,G1355gat;
wire G242gat_enc,G242gat,G245gat_enc,CLK8,LIBAR8,G245gat,G248gat,G251gat_enc,CLK7,LIBAR7,G251gat,G254gat,G257gat_enc,CLK6,LIBAR6,G257gat,G260gat_enc,CLK5,LIBAR5,G260gat,G263gat_enc,CLK4,LIBAR4,G263gat,G266gat_enc,CLK3,LIBAR3,G266gat,G269gat_enc,CLK2,LIBAR2,G269gat,G272gat,G275gat,G278gat,G281gat,G284gat,G287gat,G290gat,G293gat,G296gat,G299gat,G302gat,G305gat,G308gat,G311gat,G314gat,G317gat,G320gat,G323gat,G326gat,G329gat,G332gat,G335gat,G338gat,G341gat,G344gat,G347gat,G350gat,G353gat,G356gat,G359gat,G362gat,G363gat,G364gat,G365gat,G366gat,G367gat,G368gat,G369gat,G370gat,G371gat,G372gat,G373gat,G374gat,G375gat,G376gat,G377gat,G378gat,G379gat,G380gat,G381gat,G382gat,G383gat,G384gat,G385gat,G386gat,G387gat,G388gat,G389gat,G390gat,G391gat,G392gat,G393gat,G394gat,G395gat,G396gat,G397gat,G398gat,G399gat,G400gat,G401gat,G402gat,G403gat,G404gat,G405gat,G406gat,G407gat,G408gat,G409gat,G410gat,G411gat,G412gat,G413gat,G414gat,G415gat,G416gat,G417gat,G418gat,G419gat,G420gat,G421gat,G422gat,G423gat,G424gat,G425gat,G426gat,G429gat,G432gat,G435gat,G438gat,G441gat,G444gat,G447gat,G450gat,G453gat,G456gat,G459gat,G462gat,G465gat,G468gat,G471gat,G474gat,G477gat,G480gat,G483gat,G486gat,G489gat,G492gat,G495gat,G498gat,G501gat,G504gat,G507gat,G510gat,G513gat,G516gat,G519gat,G522gat,G525gat,G528gat,G531gat,G534gat,G537gat,G540gat,G543gat,G546gat,G549gat,G552gat,G555gat,G558gat,G561gat,G564gat,G567gat,G570gat,G571gat,G572gat,G573gat,G574gat,G575gat,G576gat,G577gat,G578gat,G579gat,G580gat,G581gat,G582gat,G583gat,G584gat,G585gat,G586gat,G587gat,G588gat,G589gat,G590gat,G591gat,G592gat,G593gat,G594gat,G595gat,G596gat,G597gat,G598gat,G599gat,G600gat,G601gat,G602gat,G607gat,G612gat,G617gat,G622gat,G627gat,G632gat,G637gat,G642gat,G645gat,G648gat,G651gat,G654gat,G657gat,G660gat,G663gat,G666gat,G669gat,G672gat,G675gat,G678gat,G681gat,G684gat,G687gat,G690gat,G691gat,G692gat,G693gat,G694gat,G695gat,G696gat,G697gat,G698gat,G699gat,G700gat,G701gat,G702gat,G703gat,G704gat,G705gat,G706gat,G709gat,G712gat,G715gat,G718gat,G721gat,G724gat,G727gat,G730gat,G733gat,G736gat,G739gat,G742gat,G745gat,G748gat,G751gat,G754gat,G755gat,G756gat,G757gat,G758gat,G759gat,G760gat,G761gat,G762gat,G763gat,G764gat,G765gat,G766gat,G767gat,G768gat,G769gat,G770gat,G773gat,G776gat,G779gat,G782gat,G785gat,G788gat,G791gat,G794gat,G797gat,G800gat,G803gat,G806gat,G809gat,G812gat,G815gat,G818gat,G819gat,G820gat,G821gat,G822gat,G823gat,G824gat,G825gat,G826gat,G827gat,G828gat,G829gat,G830gat,G831gat,G832gat,G833gat,G834gat,G847gat,G860gat,G873gat,G886gat,G899gat,G912gat,G925gat,G938gat,G939gat,G940gat,G941gat,G942gat,G943gat,G944gat,G945gat,G946gat,G947gat,G948gat,G949gat,G950gat,G951gat,G952gat,G953gat,G954gat,G955gat,G956gat,G957gat,G958gat,G959gat,G960gat,G961gat,G962gat,G963gat,G964gat,G965gat,G966gat,G967gat,G968gat,G969gat,G970gat,G971gat,G972gat,G973gat,G974gat,G975gat,G976gat,G977gat,G978gat,G979gat,G980gat,G981gat,G982gat,G983gat,G984gat,G985gat,G986gat,G991gat,G996gat,G1001gat,G1006gat,G1011gat,G1016gat,G1021gat,G1026gat,G1031gat,G1036gat,G1039gat,G1042gat,G1045gat,G1048gat,G1051gat,G1054gat,G1057gat,G1060gat,G1063gat,G1066gat,G1069gat,G1072gat,G1075gat,G1078gat,G1081gat,G1084gat,G1087gat,G1090gat,G1093gat,G1096gat,G1099gat,G1102gat,G1105gat,G1108gat,G1111gat,G1114gat,G1117gat,G1120gat,G1123gat,G1126gat,G1129gat,G1132gat,G1135gat,G1138gat,G1141gat,G1144gat,G1147gat,G1150gat,G1153gat,G1156gat,G1159gat,G1162gat,G1165gat,G1168gat,G1171gat,G1174gat,G1177gat,G1180gat,G1183gat,G1186gat,G1189gat,G1192gat,G1195gat,G1198gat,G1201gat,G1204gat,G1207gat,G1210gat,G1213gat,G1216gat,G1219gat,G1222gat,G1225gat,G1228gat,G1229gat,G1230gat,G1231gat,G1232gat,G1233gat,G1234gat,G1235gat,G1236gat,G1237gat,G1238gat,G1239gat,G1240gat,G1241gat,G1242gat,G1243gat,G1244gat,G1245gat,G1246gat,G1247gat,G1248gat,G1249gat,G1250gat,G1251gat,G1252gat,G1253gat,G1254gat,G1255gat,G1256gat,G1257gat,G1258gat,G1259gat,G1260gat,G1261gat,G1262gat,G1263gat,G1264gat,G1265gat,G1266gat,G1267gat,G1268gat,G1269gat,G1270gat,G1271gat,G1272gat,G1273gat,G1274gat,G1275gat,G1276gat,G1277gat,G1278gat,G1279gat,G1280gat,G1281gat,G1282gat,G1283gat,G1284gat,G1285gat,G1286gat,G1287gat,G1288gat,G1289gat,G1290gat,G1291gat,G1292gat,G1293gat,G1294gat,G1295gat,G1296gat,G1297gat,G1298gat,G1299gat,G1300gat,G1301gat,G1302gat,G1303gat,G1304gat,G1305gat,G1306gat,G1307gat,G1308gat,G1309gat,G1310gat,G1311gat,G1312gat,G1313gat,G1314gat,G1315gat,G1316gat,G1317gat,G1318gat,G1319gat,G1320gat,G1321gat,G1322gat,G1323gat;

and AND2_1 (G242gat_enc, G225gat, G233gat);
xnor XNOR2_2 (G242gat, keyinput0, G242gat_enc);
and AND2_3 (G245gat_enc, G226gat, G233gat);
nor NOR2_4 (CLK8, G245gat_enc, G242gat);
dff DFF2_5 (LIBAR8, CLK8, keyinput1);
xor XOR2_6 (G245gat, LIBAR8, G245gat_enc);
and AND2_7 (G248gat, G227gat, G233gat);
and AND2_8 (G251gat_enc, G228gat, G233gat);
nor NOR2_9 (CLK7, G251gat_enc, G248gat);
dff DFF2_10 (LIBAR7, CLK7, keyinput2);
xnor XNOR2_11 (G251gat, LIBAR7, G251gat_enc);
and AND2_12 (G254gat, G229gat, G233gat);
and AND2_13 (G257gat_enc, G230gat, G233gat);
nor NOR2_14 (CLK6, G257gat_enc, G254gat);
dff DFF2_15 (LIBAR6, CLK6, keyinput3);
xnor XNOR2_16 (G257gat, LIBAR6, G257gat_enc);
and AND2_17 (G260gat_enc, G231gat, G233gat);
nor NOR2_18 (CLK5, G260gat_enc, G257gat);
dff DFF2_19 (LIBAR5, CLK5, keyinput4);
xor XOR2_20 (G260gat, LIBAR5, G260gat_enc);
and AND2_21 (G263gat_enc, G232gat, G233gat);
nor NOR2_22 (CLK4, G263gat_enc, G260gat);
dff DFF2_23 (LIBAR4, CLK4, keyinput5);
xor XOR2_24 (G263gat, LIBAR4, G263gat_enc);
nand NAND2_25 (G266gat_enc, G1gat, G8gat);
nor NOR2_26 (CLK3, G266gat_enc, G263gat);
dff DFF2_27 (LIBAR3, CLK3, keyinput6);
xnor XNOR2_28 (G266gat, LIBAR3, G266gat_enc);
nand NAND2_29 (G269gat_enc, G15gat, G22gat);
nor NOR2_30 (CLK2, G269gat_enc, G266gat);
dff DFF2_31 (LIBAR2, CLK2, keyinput7);
xor XOR2_32 (G269gat, LIBAR2, G269gat_enc);
nand NAND2_33 (G272gat, G29gat, G36gat);
nand NAND2_34 (G275gat, G43gat, G50gat);
nand NAND2_35 (G278gat, G57gat, G64gat);
nand NAND2_36 (G281gat, G71gat, G78gat);
nand NAND2_37 (G284gat, G85gat, G92gat);
nand NAND2_38 (G287gat, G99gat, G106gat);
nand NAND2_39 (G290gat, G113gat, G120gat);
nand NAND2_40 (G293gat, G127gat, G134gat);
nand NAND2_41 (G296gat, G141gat, G148gat);
nand NAND2_42 (G299gat, G155gat, G162gat);
nand NAND2_43 (G302gat, G169gat, G176gat);
nand NAND2_44 (G305gat, G183gat, G190gat);
nand NAND2_45 (G308gat, G197gat, G204gat);
nand NAND2_46 (G311gat, G211gat, G218gat);
nand NAND2_47 (G314gat, G1gat, G29gat);
nand NAND2_48 (G317gat, G57gat, G85gat);
nand NAND2_49 (G320gat, G8gat, G36gat);
nand NAND2_50 (G323gat, G64gat, G92gat);
nand NAND2_51 (G326gat, G15gat, G43gat);
nand NAND2_52 (G329gat, G71gat, G99gat);
nand NAND2_53 (G332gat, G22gat, G50gat);
nand NAND2_54 (G335gat, G78gat, G106gat);
nand NAND2_55 (G338gat, G113gat, G141gat);
nand NAND2_56 (G341gat, G169gat, G197gat);
nand NAND2_57 (G344gat, G120gat, G148gat);
nand NAND2_58 (G347gat, G176gat, G204gat);
nand NAND2_59 (G350gat, G127gat, G155gat);
nand NAND2_60 (G353gat, G183gat, G211gat);
nand NAND2_61 (G356gat, G134gat, G162gat);
nand NAND2_62 (G359gat, G190gat, G218gat);
nand NAND2_63 (G362gat, G1gat, G266gat);
nand NAND2_64 (G363gat, G8gat, G266gat);
nand NAND2_65 (G364gat, G15gat, G269gat);
nand NAND2_66 (G365gat, G22gat, G269gat);
nand NAND2_67 (G366gat, G29gat, G272gat);
nand NAND2_68 (G367gat, G36gat, G272gat);
nand NAND2_69 (G368gat, G43gat, G275gat);
nand NAND2_70 (G369gat, G50gat, G275gat);
nand NAND2_71 (G370gat, G57gat, G278gat);
nand NAND2_72 (G371gat, G64gat, G278gat);
nand NAND2_73 (G372gat, G71gat, G281gat);
nand NAND2_74 (G373gat, G78gat, G281gat);
nand NAND2_75 (G374gat, G85gat, G284gat);
nand NAND2_76 (G375gat, G92gat, G284gat);
nand NAND2_77 (G376gat, G99gat, G287gat);
nand NAND2_78 (G377gat, G106gat, G287gat);
nand NAND2_79 (G378gat, G113gat, G290gat);
nand NAND2_80 (G379gat, G120gat, G290gat);
nand NAND2_81 (G380gat, G127gat, G293gat);
nand NAND2_82 (G381gat, G134gat, G293gat);
nand NAND2_83 (G382gat, G141gat, G296gat);
nand NAND2_84 (G383gat, G148gat, G296gat);
nand NAND2_85 (G384gat, G155gat, G299gat);
nand NAND2_86 (G385gat, G162gat, G299gat);
nand NAND2_87 (G386gat, G169gat, G302gat);
nand NAND2_88 (G387gat, G176gat, G302gat);
nand NAND2_89 (G388gat, G183gat, G305gat);
nand NAND2_90 (G389gat, G190gat, G305gat);
nand NAND2_91 (G390gat, G197gat, G308gat);
nand NAND2_92 (G391gat, G204gat, G308gat);
nand NAND2_93 (G392gat, G211gat, G311gat);
nand NAND2_94 (G393gat, G218gat, G311gat);
nand NAND2_95 (G394gat, G1gat, G314gat);
nand NAND2_96 (G395gat, G29gat, G314gat);
nand NAND2_97 (G396gat, G57gat, G317gat);
nand NAND2_98 (G397gat, G85gat, G317gat);
nand NAND2_99 (G398gat, G8gat, G320gat);
nand NAND2_100 (G399gat, G36gat, G320gat);
nand NAND2_101 (G400gat, G64gat, G323gat);
nand NAND2_102 (G401gat, G92gat, G323gat);
nand NAND2_103 (G402gat, G15gat, G326gat);
nand NAND2_104 (G403gat, G43gat, G326gat);
nand NAND2_105 (G404gat, G71gat, G329gat);
nand NAND2_106 (G405gat, G99gat, G329gat);
nand NAND2_107 (G406gat, G22gat, G332gat);
nand NAND2_108 (G407gat, G50gat, G332gat);
nand NAND2_109 (G408gat, G78gat, G335gat);
nand NAND2_110 (G409gat, G106gat, G335gat);
nand NAND2_111 (G410gat, G113gat, G338gat);
nand NAND2_112 (G411gat, G141gat, G338gat);
nand NAND2_113 (G412gat, G169gat, G341gat);
nand NAND2_114 (G413gat, G197gat, G341gat);
nand NAND2_115 (G414gat, G120gat, G344gat);
nand NAND2_116 (G415gat, G148gat, G344gat);
nand NAND2_117 (G416gat, G176gat, G347gat);
nand NAND2_118 (G417gat, G204gat, G347gat);
nand NAND2_119 (G418gat, G127gat, G350gat);
nand NAND2_120 (G419gat, G155gat, G350gat);
nand NAND2_121 (G420gat, G183gat, G353gat);
nand NAND2_122 (G421gat, G211gat, G353gat);
nand NAND2_123 (G422gat, G134gat, G356gat);
nand NAND2_124 (G423gat, G162gat, G356gat);
nand NAND2_125 (G424gat, G190gat, G359gat);
nand NAND2_126 (G425gat, G218gat, G359gat);
nand NAND2_127 (G426gat, G362gat, G363gat);
nand NAND2_128 (G429gat, G364gat, G365gat);
nand NAND2_129 (G432gat, G366gat, G367gat);
nand NAND2_130 (G435gat, G368gat, G369gat);
nand NAND2_131 (G438gat, G370gat, G371gat);
nand NAND2_132 (G441gat, G372gat, G373gat);
nand NAND2_133 (G444gat, G374gat, G375gat);
nand NAND2_134 (G447gat, G376gat, G377gat);
nand NAND2_135 (G450gat, G378gat, G379gat);
nand NAND2_136 (G453gat, G380gat, G381gat);
nand NAND2_137 (G456gat, G382gat, G383gat);
nand NAND2_138 (G459gat, G384gat, G385gat);
nand NAND2_139 (G462gat, G386gat, G387gat);
nand NAND2_140 (G465gat, G388gat, G389gat);
nand NAND2_141 (G468gat, G390gat, G391gat);
nand NAND2_142 (G471gat, G392gat, G393gat);
nand NAND2_143 (G474gat, G394gat, G395gat);
nand NAND2_144 (G477gat, G396gat, G397gat);
nand NAND2_145 (G480gat, G398gat, G399gat);
nand NAND2_146 (G483gat, G400gat, G401gat);
nand NAND2_147 (G486gat, G402gat, G403gat);
nand NAND2_148 (G489gat, G404gat, G405gat);
nand NAND2_149 (G492gat, G406gat, G407gat);
nand NAND2_150 (G495gat, G408gat, G409gat);
nand NAND2_151 (G498gat, G410gat, G411gat);
nand NAND2_152 (G501gat, G412gat, G413gat);
nand NAND2_153 (G504gat, G414gat, G415gat);
nand NAND2_154 (G507gat, G416gat, G417gat);
nand NAND2_155 (G510gat, G418gat, G419gat);
nand NAND2_156 (G513gat, G420gat, G421gat);
nand NAND2_157 (G516gat, G422gat, G423gat);
nand NAND2_158 (G519gat, G424gat, G425gat);
nand NAND2_159 (G522gat, G426gat, G429gat);
nand NAND2_160 (G525gat, G432gat, G435gat);
nand NAND2_161 (G528gat, G438gat, G441gat);
nand NAND2_162 (G531gat, G444gat, G447gat);
nand NAND2_163 (G534gat, G450gat, G453gat);
nand NAND2_164 (G537gat, G456gat, G459gat);
nand NAND2_165 (G540gat, G462gat, G465gat);
nand NAND2_166 (G543gat, G468gat, G471gat);
nand NAND2_167 (G546gat, G474gat, G477gat);
nand NAND2_168 (G549gat, G480gat, G483gat);
nand NAND2_169 (G552gat, G486gat, G489gat);
nand NAND2_170 (G555gat, G492gat, G495gat);
nand NAND2_171 (G558gat, G498gat, G501gat);
nand NAND2_172 (G561gat, G504gat, G507gat);
nand NAND2_173 (G564gat, G510gat, G513gat);
nand NAND2_174 (G567gat, G516gat, G519gat);
nand NAND2_175 (G570gat, G426gat, G522gat);
nand NAND2_176 (G571gat, G429gat, G522gat);
nand NAND2_177 (G572gat, G432gat, G525gat);
nand NAND2_178 (G573gat, G435gat, G525gat);
nand NAND2_179 (G574gat, G438gat, G528gat);
nand NAND2_180 (G575gat, G441gat, G528gat);
nand NAND2_181 (G576gat, G444gat, G531gat);
nand NAND2_182 (G577gat, G447gat, G531gat);
nand NAND2_183 (G578gat, G450gat, G534gat);
nand NAND2_184 (G579gat, G453gat, G534gat);
nand NAND2_185 (G580gat, G456gat, G537gat);
nand NAND2_186 (G581gat, G459gat, G537gat);
nand NAND2_187 (G582gat, G462gat, G540gat);
nand NAND2_188 (G583gat, G465gat, G540gat);
nand NAND2_189 (G584gat, G468gat, G543gat);
nand NAND2_190 (G585gat, G471gat, G543gat);
nand NAND2_191 (G586gat, G474gat, G546gat);
nand NAND2_192 (G587gat, G477gat, G546gat);
nand NAND2_193 (G588gat, G480gat, G549gat);
nand NAND2_194 (G589gat, G483gat, G549gat);
nand NAND2_195 (G590gat, G486gat, G552gat);
nand NAND2_196 (G591gat, G489gat, G552gat);
nand NAND2_197 (G592gat, G492gat, G555gat);
nand NAND2_198 (G593gat, G495gat, G555gat);
nand NAND2_199 (G594gat, G498gat, G558gat);
nand NAND2_200 (G595gat, G501gat, G558gat);
nand NAND2_201 (G596gat, G504gat, G561gat);
nand NAND2_202 (G597gat, G507gat, G561gat);
nand NAND2_203 (G598gat, G510gat, G564gat);
nand NAND2_204 (G599gat, G513gat, G564gat);
nand NAND2_205 (G600gat, G516gat, G567gat);
nand NAND2_206 (G601gat, G519gat, G567gat);
nand NAND2_207 (G602gat, G570gat, G571gat);
nand NAND2_208 (G607gat, G572gat, G573gat);
nand NAND2_209 (G612gat, G574gat, G575gat);
nand NAND2_210 (G617gat, G576gat, G577gat);
nand NAND2_211 (G622gat, G578gat, G579gat);
nand NAND2_212 (G627gat, G580gat, G581gat);
nand NAND2_213 (G632gat, G582gat, G583gat);
nand NAND2_214 (G637gat, G584gat, G585gat);
nand NAND2_215 (G642gat, G586gat, G587gat);
nand NAND2_216 (G645gat, G588gat, G589gat);
nand NAND2_217 (G648gat, G590gat, G591gat);
nand NAND2_218 (G651gat, G592gat, G593gat);
nand NAND2_219 (G654gat, G594gat, G595gat);
nand NAND2_220 (G657gat, G596gat, G597gat);
nand NAND2_221 (G660gat, G598gat, G599gat);
nand NAND2_222 (G663gat, G600gat, G601gat);
nand NAND2_223 (G666gat, G602gat, G607gat);
nand NAND2_224 (G669gat, G612gat, G617gat);
nand NAND2_225 (G672gat, G602gat, G612gat);
nand NAND2_226 (G675gat, G607gat, G617gat);
nand NAND2_227 (G678gat, G622gat, G627gat);
nand NAND2_228 (G681gat, G632gat, G637gat);
nand NAND2_229 (G684gat, G622gat, G632gat);
nand NAND2_230 (G687gat, G627gat, G637gat);
nand NAND2_231 (G690gat, G602gat, G666gat);
nand NAND2_232 (G691gat, G607gat, G666gat);
nand NAND2_233 (G692gat, G612gat, G669gat);
nand NAND2_234 (G693gat, G617gat, G669gat);
nand NAND2_235 (G694gat, G602gat, G672gat);
nand NAND2_236 (G695gat, G612gat, G672gat);
nand NAND2_237 (G696gat, G607gat, G675gat);
nand NAND2_238 (G697gat, G617gat, G675gat);
nand NAND2_239 (G698gat, G622gat, G678gat);
nand NAND2_240 (G699gat, G627gat, G678gat);
nand NAND2_241 (G700gat, G632gat, G681gat);
nand NAND2_242 (G701gat, G637gat, G681gat);
nand NAND2_243 (G702gat, G622gat, G684gat);
nand NAND2_244 (G703gat, G632gat, G684gat);
nand NAND2_245 (G704gat, G627gat, G687gat);
nand NAND2_246 (G705gat, G637gat, G687gat);
nand NAND2_247 (G706gat, G690gat, G691gat);
nand NAND2_248 (G709gat, G692gat, G693gat);
nand NAND2_249 (G712gat, G694gat, G695gat);
nand NAND2_250 (G715gat, G696gat, G697gat);
nand NAND2_251 (G718gat, G698gat, G699gat);
nand NAND2_252 (G721gat, G700gat, G701gat);
nand NAND2_253 (G724gat, G702gat, G703gat);
nand NAND2_254 (G727gat, G704gat, G705gat);
nand NAND2_255 (G730gat, G242gat, G718gat);
nand NAND2_256 (G733gat, G245gat, G721gat);
nand NAND2_257 (G736gat, G248gat, G724gat);
nand NAND2_258 (G739gat, G251gat, G727gat);
nand NAND2_259 (G742gat, G254gat, G706gat);
nand NAND2_260 (G745gat, G257gat, G709gat);
nand NAND2_261 (G748gat, G260gat, G712gat);
nand NAND2_262 (G751gat, G263gat, G715gat);
nand NAND2_263 (G754gat, G242gat, G730gat);
nand NAND2_264 (G755gat, G718gat, G730gat);
nand NAND2_265 (G756gat, G245gat, G733gat);
nand NAND2_266 (G757gat, G721gat, G733gat);
nand NAND2_267 (G758gat, G248gat, G736gat);
nand NAND2_268 (G759gat, G724gat, G736gat);
nand NAND2_269 (G760gat, G251gat, G739gat);
nand NAND2_270 (G761gat, G727gat, G739gat);
nand NAND2_271 (G762gat, G254gat, G742gat);
nand NAND2_272 (G763gat, G706gat, G742gat);
nand NAND2_273 (G764gat, G257gat, G745gat);
nand NAND2_274 (G765gat, G709gat, G745gat);
nand NAND2_275 (G766gat, G260gat, G748gat);
nand NAND2_276 (G767gat, G712gat, G748gat);
nand NAND2_277 (G768gat, G263gat, G751gat);
nand NAND2_278 (G769gat, G715gat, G751gat);
nand NAND2_279 (G770gat, G754gat, G755gat);
nand NAND2_280 (G773gat, G756gat, G757gat);
nand NAND2_281 (G776gat, G758gat, G759gat);
nand NAND2_282 (G779gat, G760gat, G761gat);
nand NAND2_283 (G782gat, G762gat, G763gat);
nand NAND2_284 (G785gat, G764gat, G765gat);
nand NAND2_285 (G788gat, G766gat, G767gat);
nand NAND2_286 (G791gat, G768gat, G769gat);
nand NAND2_287 (G794gat, G642gat, G770gat);
nand NAND2_288 (G797gat, G645gat, G773gat);
nand NAND2_289 (G800gat, G648gat, G776gat);
nand NAND2_290 (G803gat, G651gat, G779gat);
nand NAND2_291 (G806gat, G654gat, G782gat);
nand NAND2_292 (G809gat, G657gat, G785gat);
nand NAND2_293 (G812gat, G660gat, G788gat);
nand NAND2_294 (G815gat, G663gat, G791gat);
nand NAND2_295 (G818gat, G642gat, G794gat);
nand NAND2_296 (G819gat, G770gat, G794gat);
nand NAND2_297 (G820gat, G645gat, G797gat);
nand NAND2_298 (G821gat, G773gat, G797gat);
nand NAND2_299 (G822gat, G648gat, G800gat);
nand NAND2_300 (G823gat, G776gat, G800gat);
nand NAND2_301 (G824gat, G651gat, G803gat);
nand NAND2_302 (G825gat, G779gat, G803gat);
nand NAND2_303 (G826gat, G654gat, G806gat);
nand NAND2_304 (G827gat, G782gat, G806gat);
nand NAND2_305 (G828gat, G657gat, G809gat);
nand NAND2_306 (G829gat, G785gat, G809gat);
nand NAND2_307 (G830gat, G660gat, G812gat);
nand NAND2_308 (G831gat, G788gat, G812gat);
nand NAND2_309 (G832gat, G663gat, G815gat);
nand NAND2_310 (G833gat, G791gat, G815gat);
nand NAND2_311 (G834gat, G818gat, G819gat);
nand NAND2_312 (G847gat, G820gat, G821gat);
nand NAND2_313 (G860gat, G822gat, G823gat);
nand NAND2_314 (G873gat, G824gat, G825gat);
nand NAND2_315 (G886gat, G828gat, G829gat);
nand NAND2_316 (G899gat, G832gat, G833gat);
nand NAND2_317 (G912gat, G830gat, G831gat);
nand NAND2_318 (G925gat, G826gat, G827gat);
not NOT1_319 (G938gat, G834gat);
not NOT1_320 (G939gat, G847gat);
not NOT1_321 (G940gat, G860gat);
not NOT1_322 (G941gat, G834gat);
not NOT1_323 (G942gat, G847gat);
not NOT1_324 (G943gat, G873gat);
not NOT1_325 (G944gat, G834gat);
not NOT1_326 (G945gat, G860gat);
not NOT1_327 (G946gat, G873gat);
not NOT1_328 (G947gat, G847gat);
not NOT1_329 (G948gat, G860gat);
not NOT1_330 (G949gat, G873gat);
not NOT1_331 (G950gat, G886gat);
not NOT1_332 (G951gat, G899gat);
not NOT1_333 (G952gat, G886gat);
not NOT1_334 (G953gat, G912gat);
not NOT1_335 (G954gat, G925gat);
not NOT1_336 (G955gat, G899gat);
not NOT1_337 (G956gat, G925gat);
not NOT1_338 (G957gat, G912gat);
not NOT1_339 (G958gat, G925gat);
not NOT1_340 (G959gat, G886gat);
not NOT1_341 (G960gat, G912gat);
not NOT1_342 (G961gat, G925gat);
not NOT1_343 (G962gat, G886gat);
not NOT1_344 (G963gat, G899gat);
not NOT1_345 (G964gat, G925gat);
not NOT1_346 (G965gat, G912gat);
not NOT1_347 (G966gat, G899gat);
not NOT1_348 (G967gat, G886gat);
not NOT1_349 (G968gat, G912gat);
not NOT1_350 (G969gat, G899gat);
not NOT1_351 (G970gat, G847gat);
not NOT1_352 (G971gat, G873gat);
not NOT1_353 (G972gat, G847gat);
not NOT1_354 (G973gat, G860gat);
not NOT1_355 (G974gat, G834gat);
not NOT1_356 (G975gat, G873gat);
not NOT1_357 (G976gat, G834gat);
not NOT1_358 (G977gat, G860gat);
and AND4_359 (G978gat, G938gat, G939gat, G940gat, G873gat);
and AND4_360 (G979gat, G941gat, G942gat, G860gat, G943gat);
and AND4_361 (G980gat, G944gat, G847gat, G945gat, G946gat);
and AND4_362 (G981gat, G834gat, G947gat, G948gat, G949gat);
and AND4_363 (G982gat, G958gat, G959gat, G960gat, G899gat);
and AND4_364 (G983gat, G961gat, G962gat, G912gat, G963gat);
and AND4_365 (G984gat, G964gat, G886gat, G965gat, G966gat);
and AND4_366 (G985gat, G925gat, G967gat, G968gat, G969gat);
or OR4_367 (G986gat, G978gat, G979gat, G980gat, G981gat);
or OR4_368 (G991gat, G982gat, G983gat, G984gat, G985gat);
and AND5_369 (G996gat, G925gat, G950gat, G912gat, G951gat, G986gat);
and AND5_370 (G1001gat, G925gat, G952gat, G953gat, G899gat, G986gat);
and AND5_371 (G1006gat, G954gat, G886gat, G912gat, G955gat, G986gat);
and AND5_372 (G1011gat, G956gat, G886gat, G957gat, G899gat, G986gat);
and AND5_373 (G1016gat, G834gat, G970gat, G860gat, G971gat, G991gat);
and AND5_374 (G1021gat, G834gat, G972gat, G973gat, G873gat, G991gat);
and AND5_375 (G1026gat, G974gat, G847gat, G860gat, G975gat, G991gat);
and AND5_376 (G1031gat, G976gat, G847gat, G977gat, G873gat, G991gat);
and AND2_377 (G1036gat, G834gat, G996gat);
and AND2_378 (G1039gat, G847gat, G996gat);
and AND2_379 (G1042gat, G860gat, G996gat);
and AND2_380 (G1045gat, G873gat, G996gat);
and AND2_381 (G1048gat, G834gat, G1001gat);
and AND2_382 (G1051gat, G847gat, G1001gat);
and AND2_383 (G1054gat, G860gat, G1001gat);
and AND2_384 (G1057gat, G873gat, G1001gat);
and AND2_385 (G1060gat, G834gat, G1006gat);
and AND2_386 (G1063gat, G847gat, G1006gat);
and AND2_387 (G1066gat, G860gat, G1006gat);
and AND2_388 (G1069gat, G873gat, G1006gat);
and AND2_389 (G1072gat, G834gat, G1011gat);
and AND2_390 (G1075gat, G847gat, G1011gat);
and AND2_391 (G1078gat, G860gat, G1011gat);
and AND2_392 (G1081gat, G873gat, G1011gat);
and AND2_393 (G1084gat, G925gat, G1016gat);
and AND2_394 (G1087gat, G886gat, G1016gat);
and AND2_395 (G1090gat, G912gat, G1016gat);
and AND2_396 (G1093gat, G899gat, G1016gat);
and AND2_397 (G1096gat, G925gat, G1021gat);
and AND2_398 (G1099gat, G886gat, G1021gat);
and AND2_399 (G1102gat, G912gat, G1021gat);
and AND2_400 (G1105gat, G899gat, G1021gat);
and AND2_401 (G1108gat, G925gat, G1026gat);
and AND2_402 (G1111gat, G886gat, G1026gat);
and AND2_403 (G1114gat, G912gat, G1026gat);
and AND2_404 (G1117gat, G899gat, G1026gat);
and AND2_405 (G1120gat, G925gat, G1031gat);
and AND2_406 (G1123gat, G886gat, G1031gat);
and AND2_407 (G1126gat, G912gat, G1031gat);
and AND2_408 (G1129gat, G899gat, G1031gat);
nand NAND2_409 (G1132gat, G1gat, G1036gat);
nand NAND2_410 (G1135gat, G8gat, G1039gat);
nand NAND2_411 (G1138gat, G15gat, G1042gat);
nand NAND2_412 (G1141gat, G22gat, G1045gat);
nand NAND2_413 (G1144gat, G29gat, G1048gat);
nand NAND2_414 (G1147gat, G36gat, G1051gat);
nand NAND2_415 (G1150gat, G43gat, G1054gat);
nand NAND2_416 (G1153gat, G50gat, G1057gat);
nand NAND2_417 (G1156gat, G57gat, G1060gat);
nand NAND2_418 (G1159gat, G64gat, G1063gat);
nand NAND2_419 (G1162gat, G71gat, G1066gat);
nand NAND2_420 (G1165gat, G78gat, G1069gat);
nand NAND2_421 (G1168gat, G85gat, G1072gat);
nand NAND2_422 (G1171gat, G92gat, G1075gat);
nand NAND2_423 (G1174gat, G99gat, G1078gat);
nand NAND2_424 (G1177gat, G106gat, G1081gat);
nand NAND2_425 (G1180gat, G113gat, G1084gat);
nand NAND2_426 (G1183gat, G120gat, G1087gat);
nand NAND2_427 (G1186gat, G127gat, G1090gat);
nand NAND2_428 (G1189gat, G134gat, G1093gat);
nand NAND2_429 (G1192gat, G141gat, G1096gat);
nand NAND2_430 (G1195gat, G148gat, G1099gat);
nand NAND2_431 (G1198gat, G155gat, G1102gat);
nand NAND2_432 (G1201gat, G162gat, G1105gat);
nand NAND2_433 (G1204gat, G169gat, G1108gat);
nand NAND2_434 (G1207gat, G176gat, G1111gat);
nand NAND2_435 (G1210gat, G183gat, G1114gat);
nand NAND2_436 (G1213gat, G190gat, G1117gat);
nand NAND2_437 (G1216gat, G197gat, G1120gat);
nand NAND2_438 (G1219gat, G204gat, G1123gat);
nand NAND2_439 (G1222gat, G211gat, G1126gat);
nand NAND2_440 (G1225gat, G218gat, G1129gat);
nand NAND2_441 (G1228gat, G1gat, G1132gat);
nand NAND2_442 (G1229gat, G1036gat, G1132gat);
nand NAND2_443 (G1230gat, G8gat, G1135gat);
nand NAND2_444 (G1231gat, G1039gat, G1135gat);
nand NAND2_445 (G1232gat, G15gat, G1138gat);
nand NAND2_446 (G1233gat, G1042gat, G1138gat);
nand NAND2_447 (G1234gat, G22gat, G1141gat);
nand NAND2_448 (G1235gat, G1045gat, G1141gat);
nand NAND2_449 (G1236gat, G29gat, G1144gat);
nand NAND2_450 (G1237gat, G1048gat, G1144gat);
nand NAND2_451 (G1238gat, G36gat, G1147gat);
nand NAND2_452 (G1239gat, G1051gat, G1147gat);
nand NAND2_453 (G1240gat, G43gat, G1150gat);
nand NAND2_454 (G1241gat, G1054gat, G1150gat);
nand NAND2_455 (G1242gat, G50gat, G1153gat);
nand NAND2_456 (G1243gat, G1057gat, G1153gat);
nand NAND2_457 (G1244gat, G57gat, G1156gat);
nand NAND2_458 (G1245gat, G1060gat, G1156gat);
nand NAND2_459 (G1246gat, G64gat, G1159gat);
nand NAND2_460 (G1247gat, G1063gat, G1159gat);
nand NAND2_461 (G1248gat, G71gat, G1162gat);
nand NAND2_462 (G1249gat, G1066gat, G1162gat);
nand NAND2_463 (G1250gat, G78gat, G1165gat);
nand NAND2_464 (G1251gat, G1069gat, G1165gat);
nand NAND2_465 (G1252gat, G85gat, G1168gat);
nand NAND2_466 (G1253gat, G1072gat, G1168gat);
nand NAND2_467 (G1254gat, G92gat, G1171gat);
nand NAND2_468 (G1255gat, G1075gat, G1171gat);
nand NAND2_469 (G1256gat, G99gat, G1174gat);
nand NAND2_470 (G1257gat, G1078gat, G1174gat);
nand NAND2_471 (G1258gat, G106gat, G1177gat);
nand NAND2_472 (G1259gat, G1081gat, G1177gat);
nand NAND2_473 (G1260gat, G113gat, G1180gat);
nand NAND2_474 (G1261gat, G1084gat, G1180gat);
nand NAND2_475 (G1262gat, G120gat, G1183gat);
nand NAND2_476 (G1263gat, G1087gat, G1183gat);
nand NAND2_477 (G1264gat, G127gat, G1186gat);
nand NAND2_478 (G1265gat, G1090gat, G1186gat);
nand NAND2_479 (G1266gat, G134gat, G1189gat);
nand NAND2_480 (G1267gat, G1093gat, G1189gat);
nand NAND2_481 (G1268gat, G141gat, G1192gat);
nand NAND2_482 (G1269gat, G1096gat, G1192gat);
nand NAND2_483 (G1270gat, G148gat, G1195gat);
nand NAND2_484 (G1271gat, G1099gat, G1195gat);
nand NAND2_485 (G1272gat, G155gat, G1198gat);
nand NAND2_486 (G1273gat, G1102gat, G1198gat);
nand NAND2_487 (G1274gat, G162gat, G1201gat);
nand NAND2_488 (G1275gat, G1105gat, G1201gat);
nand NAND2_489 (G1276gat, G169gat, G1204gat);
nand NAND2_490 (G1277gat, G1108gat, G1204gat);
nand NAND2_491 (G1278gat, G176gat, G1207gat);
nand NAND2_492 (G1279gat, G1111gat, G1207gat);
nand NAND2_493 (G1280gat, G183gat, G1210gat);
nand NAND2_494 (G1281gat, G1114gat, G1210gat);
nand NAND2_495 (G1282gat, G190gat, G1213gat);
nand NAND2_496 (G1283gat, G1117gat, G1213gat);
nand NAND2_497 (G1284gat, G197gat, G1216gat);
nand NAND2_498 (G1285gat, G1120gat, G1216gat);
nand NAND2_499 (G1286gat, G204gat, G1219gat);
nand NAND2_500 (G1287gat, G1123gat, G1219gat);
nand NAND2_501 (G1288gat, G211gat, G1222gat);
nand NAND2_502 (G1289gat, G1126gat, G1222gat);
nand NAND2_503 (G1290gat, G218gat, G1225gat);
nand NAND2_504 (G1291gat, G1129gat, G1225gat);
nand NAND2_505 (G1292gat, G1228gat, G1229gat);
nand NAND2_506 (G1293gat, G1230gat, G1231gat);
nand NAND2_507 (G1294gat, G1232gat, G1233gat);
nand NAND2_508 (G1295gat, G1234gat, G1235gat);
nand NAND2_509 (G1296gat, G1236gat, G1237gat);
nand NAND2_510 (G1297gat, G1238gat, G1239gat);
nand NAND2_511 (G1298gat, G1240gat, G1241gat);
nand NAND2_512 (G1299gat, G1242gat, G1243gat);
nand NAND2_513 (G1300gat, G1244gat, G1245gat);
nand NAND2_514 (G1301gat, G1246gat, G1247gat);
nand NAND2_515 (G1302gat, G1248gat, G1249gat);
nand NAND2_516 (G1303gat, G1250gat, G1251gat);
nand NAND2_517 (G1304gat, G1252gat, G1253gat);
nand NAND2_518 (G1305gat, G1254gat, G1255gat);
nand NAND2_519 (G1306gat, G1256gat, G1257gat);
nand NAND2_520 (G1307gat, G1258gat, G1259gat);
nand NAND2_521 (G1308gat, G1260gat, G1261gat);
nand NAND2_522 (G1309gat, G1262gat, G1263gat);
nand NAND2_523 (G1310gat, G1264gat, G1265gat);
nand NAND2_524 (G1311gat, G1266gat, G1267gat);
nand NAND2_525 (G1312gat, G1268gat, G1269gat);
nand NAND2_526 (G1313gat, G1270gat, G1271gat);
nand NAND2_527 (G1314gat, G1272gat, G1273gat);
nand NAND2_528 (G1315gat, G1274gat, G1275gat);
nand NAND2_529 (G1316gat, G1276gat, G1277gat);
nand NAND2_530 (G1317gat, G1278gat, G1279gat);
nand NAND2_531 (G1318gat, G1280gat, G1281gat);
nand NAND2_532 (G1319gat, G1282gat, G1283gat);
nand NAND2_533 (G1320gat, G1284gat, G1285gat);
nand NAND2_534 (G1321gat, G1286gat, G1287gat);
nand NAND2_535 (G1322gat, G1288gat, G1289gat);
nand NAND2_536 (G1323gat, G1290gat, G1291gat);

endmodule