module DFF(Q, clk, D);
input D;
input clk;
output Q;
always @(clk)
begin
  Q <= D;
end
endmodule


module c432_libar_32k(G1gat,G4gat,G8gat,G11gat,G14gat,G17gat,G21gat,G24gat,G27gat,G30gat,G34gat,G37gat,G40gat,G43gat,G47gat,G50gat,G53gat,G56gat,G60gat,G63gat,G66gat,G69gat,G73gat,G76gat,G79gat,G82gat,G86gat,G89gat,G92gat,G95gat,G99gat,G102gat,G105gat,G108gat,G112gat,G115gat,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,G223gat,G329gat,G370gat,G421gat,G430gat,G431gat,G432gat);

input G1gat,G4gat,G8gat,G11gat,G14gat,G17gat,G21gat,G24gat,G27gat,G30gat,G34gat,G37gat,G40gat,G43gat,G47gat,G50gat,G53gat,G56gat,G60gat,G63gat,G66gat,G69gat,G73gat,G76gat,G79gat,G82gat,G86gat,G89gat,G92gat,G95gat,G99gat,G102gat,G105gat,G108gat,G112gat,G115gat,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31;
output G223gat,G329gat,G370gat,G421gat,G430gat,G431gat,G432gat;
wire G118gat,G119gat_enc,G119gat,G122gat_enc,CLK11,LIBAR11,G122gat,G123gat_enc,G123gat,G126gat,G127gat_enc,CLK10,LIBAR10,G127gat,G130gat,G131gat_enc,CLK9,LIBAR9,G131gat,G134gat_enc,G134gat,G135gat_enc,G135gat,G138gat_enc,G138gat,G139gat_enc,G139gat,G142gat,G143gat_enc,CLK8,LIBAR8,G143gat,G146gat_enc,CLK7,LIBAR7,G146gat,G147gat,G150gat_enc,G150gat,G151gat,G154gat,G157gat,G158gat,G159gat,G162gat_enc,CLK6,LIBAR6,G162gat,G165gat_enc,G165gat,G168gat,G171gat_enc,G171gat,G174gat_enc,CLK5,LIBAR5,G174gat,G177gat,G180gat,G183gat_enc,G183gat,G184gat_enc,G184gat,G185gat_enc,CLK4,LIBAR4,G185gat,G186gat_enc,G186gat,G187gat,G188gat,G189gat_enc,CLK3,LIBAR3,G189gat,G190gat,G191gat,G192gat,G193gat_enc,G193gat,G194gat_enc,CLK2,LIBAR2,G194gat,G195gat,G196gat,G197gat_enc,CLK1,LIBAR1,G197gat,G198gat_enc,G198gat,G1980gat,G1981gat_enc,G1981gat,G199gat_enc,G199gat,G203gat_enc,G203gat,G213gat_enc,G213gat,G224gat,G227gat_enc,G227gat,G230gat_enc,G230gat,G233gat,G236gat,G239gat,G242gat,G243gat,G246gat,G247gat,G250gat,G251gat,G254gat_enc,G254gat,G255gat,G256gat,G257gat,G258gat,G259gat,G260gat,G263gat,G264gat,G267gat,G270gat,G273gat,G276gat,G279gat,G282gat,G285gat,G288gat,G289gat,G290gat,G291gat,G292gat,G293gat,G294gat,G295gat,G2950gat,G2951gat,G296gat,G300gat,G301gat,G302gat,G303gat,G304gat,G305gat,G306gat,G307gat,G308gat,G309gat,G319gat,G330gat,G331gat,G332gat,G333gat,G334gat,G335gat,G336gat,G337gat,G338gat,G339gat,G340gat,G341gat,G342gat,G343gat,G344gat,G345gat,G346gat,G347gat,G348gat,G349gat,G350gat,G351gat,G352gat,G353gat,G354gat,G355gat,G356gat,G3560gat,G3561gat,G357gat,G360gat,G371gat,G372gat,G373gat,G374gat,G375gat,G376gat,G377gat,G378gat,G379gat,G380gat,G381gat,G386gat,G393gat,G399gat,G404gat,G407gat,G411gat,G414gat,G415gat,G4150gat,G4151gat,G416gat,G417gat,G418gat,G419gat,G420gat,G422gat,G425gat,G428gat,G429gat;

not NOT1_1 (G118gat, G1gat);
not NOT1_2 (G119gat_enc, G4gat);
xnor XNOR2_3 (G119gat, keyinput0, G119gat_enc);
not NOT1_4 (G122gat_enc, G11gat);
nor NOR2_5 (CLK11, G122gat_enc, G119gat);
dff DFF2_6 (LIBAR11, CLK11, keyinput1);
xor XOR2_7 (G122gat, LIBAR11, G122gat_enc);
not NOT1_8 (G123gat_enc, G17gat);
xor XOR2_9 (G123gat, keyinput2, G123gat_enc);
not NOT1_10 (G126gat, G24gat);
not NOT1_11 (G127gat_enc, G30gat);
nor NOR2_12 (CLK10, G127gat_enc, G126gat);
dff DFF2_13 (LIBAR10, CLK10, keyinput3);
xnor XNOR2_14 (G127gat, LIBAR10, G127gat_enc);
not NOT1_15 (G130gat, G37gat);
not NOT1_16 (G131gat_enc, G43gat);
nor NOR2_17 (CLK9, G131gat_enc, G130gat);
dff DFF2_18 (LIBAR9, CLK9, keyinput4);
xnor XNOR2_19 (G131gat, LIBAR9, G131gat_enc);
not NOT1_20 (G134gat_enc, G50gat);
xor XOR2_21 (G134gat, keyinput5, G134gat_enc);
not NOT1_22 (G135gat_enc, G56gat);
xor XOR2_23 (G135gat, keyinput6, G135gat_enc);
not NOT1_24 (G138gat_enc, G63gat);
xor XOR2_25 (G138gat, keyinput7, G138gat_enc);
not NOT1_26 (G139gat_enc, G69gat);
xnor XNOR2_27 (G139gat, keyinput8, G139gat_enc);
not NOT1_28 (G142gat, G76gat);
not NOT1_29 (G143gat_enc, G82gat);
nor NOR2_30 (CLK8, G143gat_enc, G142gat);
dff DFF2_31 (LIBAR8, CLK8, keyinput9);
xnor XNOR2_32 (G143gat, LIBAR8, G143gat_enc);
not NOT1_33 (G146gat_enc, G89gat);
nor NOR2_34 (CLK7, G146gat_enc, G143gat);
dff DFF2_35 (LIBAR7, CLK7, keyinput10);
xnor XNOR2_36 (G146gat, LIBAR7, G146gat_enc);
not NOT1_37 (G147gat, G95gat);
not NOT1_38 (G150gat_enc, G102gat);
xnor XNOR2_39 (G150gat, keyinput11, G150gat_enc);
not NOT1_40 (G151gat, G108gat);
nand NAND2_41 (G154gat, G118gat, G4gat);
nor NOR2_42 (G157gat, G8gat, G119gat);
nor NOR2_43 (G158gat, G14gat, G119gat);
nand NAND2_44 (G159gat, G122gat, G17gat);
nand NAND2_45 (G162gat_enc, G126gat, G30gat);
nor NOR2_46 (CLK6, G162gat_enc, G159gat);
dff DFF2_47 (LIBAR6, CLK6, keyinput12);
xnor XNOR2_48 (G162gat, LIBAR6, G162gat_enc);
nand NAND2_49 (G165gat_enc, G130gat, G43gat);
xor XOR2_50 (G165gat, keyinput13, G165gat_enc);
nand NAND2_51 (G168gat, G134gat, G56gat);
nand NAND2_52 (G171gat_enc, G138gat, G69gat);
xnor XNOR2_53 (G171gat, keyinput14, G171gat_enc);
nand NAND2_54 (G174gat_enc, G142gat, G82gat);
nor NOR2_55 (CLK5, G174gat_enc, G171gat);
dff DFF2_56 (LIBAR5, CLK5, keyinput15);
xor XOR2_57 (G174gat, LIBAR5, G174gat_enc);
nand NAND2_58 (G177gat, G146gat, G95gat);
nand NAND2_59 (G180gat, G150gat, G108gat);
nor NOR2_60 (G183gat_enc, G21gat, G123gat);
xnor XNOR2_61 (G183gat, keyinput16, G183gat_enc);
nor NOR2_62 (G184gat_enc, G27gat, G123gat);
xor XOR2_63 (G184gat, keyinput17, G184gat_enc);
nor NOR2_64 (G185gat_enc, G34gat, G127gat);
nor NOR2_65 (CLK4, G185gat_enc, G184gat);
dff DFF2_66 (LIBAR4, CLK4, keyinput18);
xnor XNOR2_67 (G185gat, LIBAR4, G185gat_enc);
nor NOR2_68 (G186gat_enc, G40gat, G127gat);
xor XOR2_69 (G186gat, keyinput19, G186gat_enc);
nor NOR2_70 (G187gat, G47gat, G131gat);
nor NOR2_71 (G188gat, G53gat, G131gat);
nor NOR2_72 (G189gat_enc, G60gat, G135gat);
nor NOR2_73 (CLK3, G189gat_enc, G188gat);
dff DFF2_74 (LIBAR3, CLK3, keyinput20);
xnor XNOR2_75 (G189gat, LIBAR3, G189gat_enc);
nor NOR2_76 (G190gat, G66gat, G135gat);
nor NOR2_77 (G191gat, G73gat, G139gat);
nor NOR2_78 (G192gat, G79gat, G139gat);
nor NOR2_79 (G193gat_enc, G86gat, G143gat);
xnor XNOR2_80 (G193gat, keyinput21, G193gat_enc);
nor NOR2_81 (G194gat_enc, G92gat, G143gat);
nor NOR2_82 (CLK2, G194gat_enc, G193gat);
dff DFF2_83 (LIBAR2, CLK2, keyinput22);
xnor XNOR2_84 (G194gat, LIBAR2, G194gat_enc);
nor NOR2_85 (G195gat, G99gat, G147gat);
nor NOR2_86 (G196gat, G105gat, G147gat);
nor NOR2_87 (G197gat_enc, G112gat, G151gat);
nor NOR2_88 (CLK1, G197gat_enc, G196gat);
dff DFF2_89 (LIBAR1, CLK1, keyinput23);
xnor XNOR2_90 (G197gat, LIBAR1, G197gat_enc);
nor NOR2_91 (G198gat_enc, G115gat, G151gat);
xor XOR2_92 (G198gat, keyinput24, G198gat_enc);
and AND4_93 (G1980gat, G154gat, G159gat, G162gat, G165gat);
and AND5_94 (G1981gat_enc, G168gat, G171gat, G174gat, G177gat, G180gat);
xnor XNOR2_95 (G1981gat, keyinput25, G1981gat_enc);
and AND2_96 (G199gat_enc, G1980gat, G1981gat);
xor XOR2_97 (G199gat, keyinput26, G199gat_enc);
not NOT1_98 (G203gat_enc, G199gat);
xnor XNOR2_99 (G203gat, keyinput27, G203gat_enc);
not NOT1_100 (G213gat_enc, G199gat);
xor XOR2_101 (G213gat, keyinput28, G213gat_enc);
not NOT1_102 (G223gat, G199gat);
xor XOR2_103 (G224gat, G203gat, G154gat);
xor XOR2_104 (G227gat_enc, G203gat, G159gat);
xnor XNOR2_105 (G227gat, keyinput29, G227gat_enc);
xor XOR2_106 (G230gat_enc, G203gat, G162gat);
xor XOR2_107 (G230gat, keyinput30, G230gat_enc);
xor XOR2_108 (G233gat, G203gat, G165gat);
xor XOR2_109 (G236gat, G203gat, G168gat);
xor XOR2_110 (G239gat, G203gat, G171gat);
nand NAND2_111 (G242gat, G1gat, G213gat);
xor XOR2_112 (G243gat, G203gat, G174gat);
nand NAND2_113 (G246gat, G213gat, G11gat);
xor XOR2_114 (G247gat, G203gat, G177gat);
nand NAND2_115 (G250gat, G213gat, G24gat);
xor XOR2_116 (G251gat, G203gat, G180gat);
nand NAND2_117 (G254gat_enc, G213gat, G37gat);
xnor XNOR2_118 (G254gat, keyinput31, G254gat_enc);
nand NAND2_119 (G255gat, G213gat, G50gat);
nand NAND2_120 (G256gat, G213gat, G63gat);
nand NAND2_121 (G257gat, G213gat, G76gat);
nand NAND2_122 (G258gat, G213gat, G89gat);
nand NAND2_123 (G259gat, G213gat, G102gat);
nand NAND2_124 (G260gat, G224gat, G157gat);
nand NAND2_125 (G263gat, G224gat, G158gat);
nand NAND2_126 (G264gat, G227gat, G183gat);
nand NAND2_127 (G267gat, G230gat, G185gat);
nand NAND2_128 (G270gat, G233gat, G187gat);
nand NAND2_129 (G273gat, G236gat, G189gat);
nand NAND2_130 (G276gat, G239gat, G191gat);
nand NAND2_131 (G279gat, G243gat, G193gat);
nand NAND2_132 (G282gat, G247gat, G195gat);
nand NAND2_133 (G285gat, G251gat, G197gat);
nand NAND2_134 (G288gat, G227gat, G184gat);
nand NAND2_135 (G289gat, G230gat, G186gat);
nand NAND2_136 (G290gat, G233gat, G188gat);
nand NAND2_137 (G291gat, G236gat, G190gat);
nand NAND2_138 (G292gat, G239gat, G192gat);
nand NAND2_139 (G293gat, G243gat, G194gat);
nand NAND2_140 (G294gat, G247gat, G196gat);
nand NAND2_141 (G295gat, G251gat, G198gat);
and AND4_142 (G2950gat, G260gat, G264gat, G267gat, G270gat);
and AND5_143 (G2951gat, G273gat, G276gat, G279gat, G282gat, G285gat);
and AND2_144 (G296gat, G2950gat, G2951gat);
not NOT1_145 (G300gat, G263gat);
not NOT1_146 (G301gat, G288gat);
not NOT1_147 (G302gat, G289gat);
not NOT1_148 (G303gat, G290gat);
not NOT1_149 (G304gat, G291gat);
not NOT1_150 (G305gat, G292gat);
not NOT1_151 (G306gat, G293gat);
not NOT1_152 (G307gat, G294gat);
not NOT1_153 (G308gat, G295gat);
not NOT1_154 (G309gat, G296gat);
not NOT1_155 (G319gat, G296gat);
not NOT1_156 (G329gat, G296gat);
xor XOR2_157 (G330gat, G309gat, G260gat);
xor XOR2_158 (G331gat, G309gat, G264gat);
xor XOR2_159 (G332gat, G309gat, G267gat);
xor XOR2_160 (G333gat, G309gat, G270gat);
nand NAND2_161 (G334gat, G8gat, G319gat);
xor XOR2_162 (G335gat, G309gat, G273gat);
nand NAND2_163 (G336gat, G319gat, G21gat);
xor XOR2_164 (G337gat, G309gat, G276gat);
nand NAND2_165 (G338gat, G319gat, G34gat);
xor XOR2_166 (G339gat, G309gat, G279gat);
nand NAND2_167 (G340gat, G319gat, G47gat);
xor XOR2_168 (G341gat, G309gat, G282gat);
nand NAND2_169 (G342gat, G319gat, G60gat);
xor XOR2_170 (G343gat, G309gat, G285gat);
nand NAND2_171 (G344gat, G319gat, G73gat);
nand NAND2_172 (G345gat, G319gat, G86gat);
nand NAND2_173 (G346gat, G319gat, G99gat);
nand NAND2_174 (G347gat, G319gat, G112gat);
nand NAND2_175 (G348gat, G330gat, G300gat);
nand NAND2_176 (G349gat, G331gat, G301gat);
nand NAND2_177 (G350gat, G332gat, G302gat);
nand NAND2_178 (G351gat, G333gat, G303gat);
nand NAND2_179 (G352gat, G335gat, G304gat);
nand NAND2_180 (G353gat, G337gat, G305gat);
nand NAND2_181 (G354gat, G339gat, G306gat);
nand NAND2_182 (G355gat, G341gat, G307gat);
nand NAND2_183 (G356gat, G343gat, G308gat);
and AND4_184 (G3560gat, G348gat, G349gat, G350gat, G351gat);
and AND5_185 (G3561gat, G352gat, G353gat, G354gat, G355gat, G356gat);
and AND2_186 (G357gat, G3560gat, G3561gat);
not NOT1_187 (G360gat, G357gat);
not NOT1_188 (G370gat, G357gat);
nand NAND2_189 (G371gat, G14gat, G360gat);
nand NAND2_190 (G372gat, G360gat, G27gat);
nand NAND2_191 (G373gat, G360gat, G40gat);
nand NAND2_192 (G374gat, G360gat, G53gat);
nand NAND2_193 (G375gat, G360gat, G66gat);
nand NAND2_194 (G376gat, G360gat, G79gat);
nand NAND2_195 (G377gat, G360gat, G92gat);
nand NAND2_196 (G378gat, G360gat, G105gat);
nand NAND2_197 (G379gat, G360gat, G115gat);
nand NAND4_198 (G380gat, G4gat, G242gat, G334gat, G371gat);
nand NAND4_199 (G381gat, G246gat, G336gat, G372gat, G17gat);
nand NAND4_200 (G386gat, G250gat, G338gat, G373gat, G30gat);
nand NAND4_201 (G393gat, G254gat, G340gat, G374gat, G43gat);
nand NAND4_202 (G399gat, G255gat, G342gat, G375gat, G56gat);
nand NAND4_203 (G404gat, G256gat, G344gat, G376gat, G69gat);
nand NAND4_204 (G407gat, G257gat, G345gat, G377gat, G82gat);
nand NAND4_205 (G411gat, G258gat, G346gat, G378gat, G95gat);
nand NAND4_206 (G414gat, G259gat, G347gat, G379gat, G108gat);
not NOT1_207 (G415gat, G380gat);
and AND4_208 (G4150gat, G381gat, G386gat, G393gat, G399gat);
and AND4_209 (G4151gat, G404gat, G407gat, G411gat, G414gat);
and AND2_210 (G416gat, G4150gat, G4151gat);
not NOT1_211 (G417gat, G393gat);
not NOT1_212 (G418gat, G404gat);
not NOT1_213 (G419gat, G407gat);
not NOT1_214 (G420gat, G411gat);
nor NOR2_215 (G421gat, G415gat, G416gat);
nand NAND2_216 (G422gat, G386gat, G417gat);
nand NAND4_217 (G425gat, G386gat, G393gat, G418gat, G399gat);
nand NAND3_218 (G428gat, G399gat, G393gat, G419gat);
nand NAND4_219 (G429gat, G386gat, G393gat, G407gat, G420gat);
nand NAND4_220 (G430gat, G381gat, G386gat, G422gat, G399gat);
nand NAND4_221 (G431gat, G381gat, G386gat, G425gat, G428gat);
nand NAND4_222 (G432gat, G381gat, G422gat, G425gat, G429gat);

endmodule