module cac(keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,n6123);

input keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31;
output n6123;
wire wire1669,wire1670,wire1347,wire1504,wire1505,wire1355,wire1673,wire1674,wire1343,wire1331,wire1500,wire1501,wire1413,wire1414,wire1421,wire1422,wire1365,wire1393,wire1323,wire1325,n_0,wire1335,wire1351,wire1353,wire1425,wire1426,wire1429,wire1430,wire1339,wire1389,wire1409,wire1410,wire1319,wire1385,wire1377,n_1,wire1397,wire1373,wire1375,wire1369,wire1371,wire1315,wire1327,wire1417,wire1418,wire1381,wire1671,wire1348,wire1349,wire1506,wire1356,wire1357,wire1675,wire1344,wire1345,wire1332,wire1333,wire1502,wire1415,wire1423,wire1366,wire1367,wire1394,wire1395,wire1324,wire1304,wire1305,wire1336,wire1337,wire1352,wire1427,wire1431,wire1340,wire1341,wire1390,wire1391,wire1411,wire1320,wire1321,wire1386,wire1387,wire1378,wire1379,wire1308,wire1309,wire1398,wire1399,wire1374,wire1370,wire1316,wire1317,wire1328,wire1329,wire1419,wire1382,wire1383,n_1524,wire1350,wire1507,wire1358,n_1525,wire1346,wire1334,wire1503,wire1416,wire1424,wire1368,wire1396,wire1326,wire1306,wire1338,wire1354,wire1428,wire1432,wire1342,wire1392,wire1412,wire1322,wire1388,wire1380,wire1310,wire1400,wire1376,wire1372,wire1318,wire1330,wire1420,wire1384,n_68,n_6,n_65,n_69,n_72,n_7,n_38,n_36,n_57,n_50,n_75,n_71,n_66,n_33,n_32,n_70,n_51,n_39,n_76,n_52,n_54,n_49,n_55,n_56,n_78,n_74,n_37,n_53,wire1295,wire1297,wire1300,wire1307,wire1298,wire1299,wire1311,wire1296,n_109,n_106,n_102,n_90,n_105,n_103,n_88,n_108,wire1260,wire1258,wire1259,n_124,n_126,n_125,wire1035,wire1036,wire1037,n_1412,wire89,wire90,wire91,wire92;

not NOT1_1 (wire1669, keyinput0);
and AND2_2 (wire1670, n256, keyinput0);
not NOT1_3 (wire1347, keyinput1);
or OR2_4 (wire1504, n239, keyinput2);
and AND2_5 (wire1505, n239, keyinput2);
not NOT1_6 (wire1355, keyinput3);
not NOT1_7 (wire1673, keyinput4);
and AND2_8 (wire1674, n222, keyinput4);
not NOT1_9 (wire1343, keyinput5);
not NOT1_10 (wire1331, keyinput6);
or OR2_11 (wire1500, n324, keyinput7);
and AND2_12 (wire1501, n324, keyinput7);
or OR2_13 (wire1413, n188, keyinput8);
and AND2_14 (wire1414, n188, keyinput8);
or OR2_15 (wire1421, n341, keyinput9);
and AND2_16 (wire1422, n341, keyinput9);
not NOT1_17 (wire1365, keyinput10);
not NOT1_18 (wire1393, keyinput11);
not NOT1_19 (wire1323, keyinput12);
and AND2_20 (wire1325, keyinput12, n154);
not NOT1_21 (n_0, keyinput13);
not NOT1_22 (wire1335, keyinput14);
not NOT1_23 (wire1351, keyinput15);
and AND2_24 (wire1353, keyinput15, n392);
or OR2_25 (wire1425, n120, keyinput16);
and AND2_26 (wire1426, n120, keyinput16);
or OR2_27 (wire1429, n409, keyinput17);
and AND2_28 (wire1430, n409, keyinput17);
not NOT1_29 (wire1339, keyinput18);
not NOT1_30 (wire1389, keyinput19);
or OR2_31 (wire1409, n86, keyinput20);
and AND2_32 (wire1410, n86, keyinput20);
not NOT1_33 (wire1319, keyinput21);
not NOT1_34 (wire1385, keyinput22);
not NOT1_35 (wire1377, keyinput23);
not NOT1_36 (n_1, keyinput24);
not NOT1_37 (wire1397, keyinput25);
not NOT1_38 (wire1373, keyinput26);
and AND2_39 (wire1375, keyinput26, n35);
not NOT1_40 (wire1369, keyinput27);
and AND2_41 (wire1371, keyinput27, n494);
not NOT1_42 (wire1315, keyinput28);
not NOT1_43 (wire1327, keyinput29);
or OR2_44 (wire1417, n528, keyinput30);
and AND2_45 (wire1418, n528, keyinput30);
not NOT1_46 (wire1381, keyinput31);
and AND2_47 (wire1671, wire1668, wire1669);
and AND2_48 (wire1348, wire1347, n290);
and AND2_49 (wire1349, keyinput1, n_67);
not NOT1_50 (wire1506, wire1505);
and AND2_51 (wire1356, wire1355, n307);
and AND2_52 (wire1357, keyinput3, n_25);
and AND2_53 (wire1675, wire1672, wire1673);
and AND2_54 (wire1344, wire1343, n273);
and AND2_55 (wire1345, keyinput5, n_8);
and AND2_56 (wire1332, wire1331, n205);
and AND2_57 (wire1333, keyinput6, n_17);
not NOT1_58 (wire1502, wire1501);
not NOT1_59 (wire1415, wire1414);
not NOT1_60 (wire1423, wire1422);
and AND2_61 (wire1366, wire1365, n171);
and AND2_62 (wire1367, keyinput10, n_21);
and AND2_63 (wire1394, wire1393, n358);
and AND2_64 (wire1395, keyinput11, n_28);
and AND2_65 (wire1324, wire1323, n_19);
or OR2_66 (wire1304, n375, n_0);
or OR2_67 (wire1305, n_89, keyinput13);
and AND2_68 (wire1336, wire1335, n137);
and AND2_69 (wire1337, keyinput14, n_20);
and AND2_70 (wire1352, wire1351, n_11);
not NOT1_71 (wire1427, wire1426);
not NOT1_72 (wire1431, wire1430);
and AND2_73 (wire1340, wire1339, n103);
and AND2_74 (wire1341, keyinput18, n_31);
and AND2_75 (wire1390, wire1389, n426);
and AND2_76 (wire1391, keyinput19, n_12);
not NOT1_77 (wire1411, wire1410);
and AND2_78 (wire1320, wire1319, n443);
and AND2_79 (wire1321, keyinput21, n_24);
and AND2_80 (wire1386, wire1385, n69);
and AND2_81 (wire1387, keyinput22, n_22);
and AND2_82 (wire1378, wire1377, n460);
and AND2_83 (wire1379, keyinput23, n_26);
or OR2_84 (wire1308, n52, n_1);
or OR2_85 (wire1309, n_87, keyinput24);
and AND2_86 (wire1398, wire1397, n477);
and AND2_87 (wire1399, keyinput25, n_30);
and AND2_88 (wire1374, wire1373, n_4);
and AND2_89 (wire1370, wire1369, n_16);
and AND2_90 (wire1316, wire1315, n18);
and AND2_91 (wire1317, keyinput28, n_77);
and AND2_92 (wire1328, wire1327, n511);
and AND2_93 (wire1329, keyinput29, n_73);
not NOT1_94 (wire1419, wire1418);
and AND2_95 (wire1382, wire1381, n1);
and AND2_96 (wire1383, keyinput31, n_9);
or OR2_97 (n_1524, wire1671, wire1670);
or OR2_98 (wire1350, wire1349, wire1348);
and AND2_99 (wire1507, wire1506, wire1504);
or OR2_100 (wire1358, wire1357, wire1356);
or OR2_101 (n_1525, wire1675, wire1674);
or OR2_102 (wire1346, wire1345, wire1344);
or OR2_103 (wire1334, wire1333, wire1332);
and AND2_104 (wire1503, wire1502, wire1500);
and AND2_105 (wire1416, wire1415, wire1413);
and AND2_106 (wire1424, wire1423, wire1421);
or OR2_107 (wire1368, wire1367, wire1366);
or OR2_108 (wire1396, wire1395, wire1394);
or OR2_109 (wire1326, wire1325, wire1324);
and AND2_110 (wire1306, wire1305, wire1304);
or OR2_111 (wire1338, wire1337, wire1336);
or OR2_112 (wire1354, wire1353, wire1352);
and AND2_113 (wire1428, wire1427, wire1425);
and AND2_114 (wire1432, wire1431, wire1429);
or OR2_115 (wire1342, wire1341, wire1340);
or OR2_116 (wire1392, wire1391, wire1390);
and AND2_117 (wire1412, wire1411, wire1409);
or OR2_118 (wire1322, wire1321, wire1320);
or OR2_119 (wire1388, wire1387, wire1386);
or OR2_120 (wire1380, wire1379, wire1378);
and AND2_121 (wire1310, wire1309, wire1308);
or OR2_122 (wire1400, wire1399, wire1398);
or OR2_123 (wire1376, wire1375, wire1374);
or OR2_124 (wire1372, wire1371, wire1370);
or OR2_125 (wire1318, wire1317, wire1316);
or OR2_126 (wire1330, wire1329, wire1328);
and AND2_127 (wire1420, wire1419, wire1417);
or OR2_128 (wire1384, wire1383, wire1382);
not NOT1_129 (n_68, wire1350);
not NOT1_130 (n_6, wire1507);
not NOT1_131 (n_65, wire1358);
not NOT1_132 (n_69, wire1346);
not NOT1_133 (n_72, wire1334);
not NOT1_134 (n_7, wire1503);
not NOT1_135 (n_38, wire1416);
not NOT1_136 (n_36, wire1424);
not NOT1_137 (n_57, wire1368);
not NOT1_138 (n_50, wire1396);
not NOT1_139 (n_75, wire1326);
not NOT1_140 (n_71, wire1338);
not NOT1_141 (n_66, wire1354);
not NOT1_142 (n_33, wire1428);
not NOT1_143 (n_32, wire1432);
not NOT1_144 (n_70, wire1342);
not NOT1_145 (n_51, wire1392);
not NOT1_146 (n_39, wire1412);
not NOT1_147 (n_76, wire1322);
not NOT1_148 (n_52, wire1388);
not NOT1_149 (n_54, wire1380);
not NOT1_150 (n_49, wire1400);
not NOT1_151 (n_55, wire1376);
not NOT1_152 (n_56, wire1372);
not NOT1_153 (n_78, wire1318);
not NOT1_154 (n_74, wire1330);
not NOT1_155 (n_37, wire1420);
not NOT1_156 (n_53, wire1384);
and AND4_157 (wire1295, n_1524, n_68, n_65, n_6);
and AND4_158 (wire1297, n_72, n_1525, n_69, n_7);
and AND4_159 (wire1300, n_57, n_50, n_36, n_38);
and AND2_160 (wire1307, wire1306, n_71);
and AND4_161 (wire1298, n_51, n_70, n_32, n_33);
and AND4_162 (wire1299, n_54, n_52, n_76, n_39);
and AND2_163 (wire1311, wire1310, n_49);
and AND4_164 (wire1296, n_53, n_74, n_78, n_37);
not NOT1_165 (n_109, wire1295);
not NOT1_166 (n_106, wire1297);
not NOT1_167 (n_102, wire1300);
not NOT1_168 (n_90, wire1307);
not NOT1_169 (n_105, wire1298);
not NOT1_170 (n_103, wire1299);
not NOT1_171 (n_88, wire1311);
not NOT1_172 (n_108, wire1296);
or OR4_173 (wire1260, n_108, n_109, n_103, n_105);
or OR4_174 (wire1258, n_106, n_90, n_75, n_66);
or OR4_175 (wire1259, n_102, n_88, n_56, n_55);
not NOT1_176 (n_124, wire1260);
not NOT1_177 (n_126, wire1258);
not NOT1_178 (n_125, wire1259);
and AND2_179 (wire1035, n_124, n_125);
and AND2_180 (wire1036, wire1035, n_126);
or OR2_181 (wire1037, wire1036, n_373);
not NOT1_182 (n_1412, wire1037);
or OR2_183 (wire89, n_1413, n_1412);
and AND2_184 (wire90, n_1413, n_1412);
not NOT1_185 (wire91, wire90);
and AND2_186 (wire92, wire91, wire89);
not NOT1_187 (n6123, wire92);

endmodule