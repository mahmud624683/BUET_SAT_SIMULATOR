module c432(G1gat,G4gat,G8gat,G11gat,G14gat,G17gat,G21gat,G24gat,G27gat,G30gat,G34gat,G37gat,G40gat,G43gat,G47gat,G50gat,G53gat,G56gat,G60gat,G63gat,G66gat,G69gat,G73gat,G76gat,G79gat,G82gat,G86gat,G89gat,G92gat,G95gat,G99gat,G102gat,G105gat,G108gat,G112gat,G115gat,G223gat,G329gat,G370gat,G421gat,G430gat,G431gat,G432gat);

input G1gat,G4gat,G8gat,G11gat,G14gat,G17gat,G21gat,G24gat,G27gat,G30gat,G34gat,G37gat,G40gat,G43gat,G47gat,G50gat,G53gat,G56gat,G60gat,G63gat,G66gat,G69gat,G73gat,G76gat,G79gat,G82gat,G86gat,G89gat,G92gat,G95gat,G99gat,G102gat,G105gat,G108gat,G112gat,G115gat;
output G223gat,G329gat,G370gat,G421gat,G430gat,G431gat,G432gat;
wire G118gat,G119gat,G122gat,G123gat,G126gat,G127gat,G130gat,G131gat,G134gat,G135gat,G138gat,G139gat,G142gat,G143gat,G146gat,G147gat,G150gat,G151gat,G154gat,G157gat,G158gat,G159gat,G162gat,G165gat,G168gat,G171gat,G174gat,G177gat,G180gat,G183gat,G184gat,G185gat,G186gat,G187gat,G188gat,G189gat,G190gat,G191gat,G192gat,G193gat,G194gat,G195gat,G196gat,G197gat,G198gat,G1980gat,G1981gat,G199gat,G203gat,G213gat,G224gat,G227gat,G230gat,G233gat,G236gat,G239gat,G242gat,G243gat,G246gat,G247gat,G250gat,G251gat,G254gat,G255gat,G256gat,G257gat,G258gat,G259gat,G260gat,G263gat,G264gat,G267gat,G270gat,G273gat,G276gat,G279gat,G282gat,G285gat,G288gat,G289gat,G290gat,G291gat,G292gat,G293gat,G294gat,G295gat,G2950gat,G2951gat,G296gat,G300gat,G301gat,G302gat,G303gat,G304gat,G305gat,G306gat,G307gat,G308gat,G309gat,G319gat,G330gat,G331gat,G332gat,G333gat,G334gat,G335gat,G336gat,G337gat,G338gat,G339gat,G340gat,G341gat,G342gat,G343gat,G344gat,G345gat,G346gat,G347gat,G348gat,G349gat,G350gat,G351gat,G352gat,G353gat,G354gat,G355gat,G356gat,G3560gat,G3561gat,G357gat,G360gat,G371gat,G372gat,G373gat,G374gat,G375gat,G376gat,G377gat,G378gat,G379gat,G380gat,G381gat,G386gat,G393gat,G399gat,G404gat,G407gat,G411gat,G414gat,G415gat,G4150gat,G4151gat,G416gat,G417gat,G418gat,G419gat,G420gat,G422gat,G425gat,G428gat,G429gat;

not NOT1_1 (G118gat, G1gat);
not NOT1_2 (G119gat, G4gat);
not NOT1_3 (G122gat, G11gat);
not NOT1_4 (G123gat, G17gat);
not NOT1_5 (G126gat, G24gat);
not NOT1_6 (G127gat, G30gat);
not NOT1_7 (G130gat, G37gat);
not NOT1_8 (G131gat, G43gat);
not NOT1_9 (G134gat, G50gat);
not NOT1_10 (G135gat, G56gat);
not NOT1_11 (G138gat, G63gat);
not NOT1_12 (G139gat, G69gat);
not NOT1_13 (G142gat, G76gat);
not NOT1_14 (G143gat, G82gat);
not NOT1_15 (G146gat, G89gat);
not NOT1_16 (G147gat, G95gat);
not NOT1_17 (G150gat, G102gat);
not NOT1_18 (G151gat, G108gat);
nand NAND2_19 (G154gat, G118gat, G4gat);
nor NOR2_20 (G157gat, G8gat, G119gat);
nor NOR2_21 (G158gat, G14gat, G119gat);
nand NAND2_22 (G159gat, G122gat, G17gat);
nand NAND2_23 (G162gat, G126gat, G30gat);
nand NAND2_24 (G165gat, G130gat, G43gat);
nand NAND2_25 (G168gat, G134gat, G56gat);
nand NAND2_26 (G171gat, G138gat, G69gat);
nand NAND2_27 (G174gat, G142gat, G82gat);
nand NAND2_28 (G177gat, G146gat, G95gat);
nand NAND2_29 (G180gat, G150gat, G108gat);
nor NOR2_30 (G183gat, G21gat, G123gat);
nor NOR2_31 (G184gat, G27gat, G123gat);
nor NOR2_32 (G185gat, G34gat, G127gat);
nor NOR2_33 (G186gat, G40gat, G127gat);
nor NOR2_34 (G187gat, G47gat, G131gat);
nor NOR2_35 (G188gat, G53gat, G131gat);
nor NOR2_36 (G189gat, G60gat, G135gat);
nor NOR2_37 (G190gat, G66gat, G135gat);
nor NOR2_38 (G191gat, G73gat, G139gat);
nor NOR2_39 (G192gat, G79gat, G139gat);
nor NOR2_40 (G193gat, G86gat, G143gat);
nor NOR2_41 (G194gat, G92gat, G143gat);
nor NOR2_42 (G195gat, G99gat, G147gat);
nor NOR2_43 (G196gat, G105gat, G147gat);
nor NOR2_44 (G197gat, G112gat, G151gat);
nor NOR2_45 (G198gat, G115gat, G151gat);
and AND4_46 (G1980gat, G154gat, G159gat, G162gat, G165gat);
and AND5_47 (G1981gat, G168gat, G171gat, G174gat, G177gat, G180gat);
and AND2_48 (G199gat, G1980gat, G1981gat);
not NOT1_49 (G203gat, G199gat);
not NOT1_50 (G213gat, G199gat);
not NOT1_51 (G223gat, G199gat);
xor XOR2_52 (G224gat, G203gat, G154gat);
xor XOR2_53 (G227gat, G203gat, G159gat);
xor XOR2_54 (G230gat, G203gat, G162gat);
xor XOR2_55 (G233gat, G203gat, G165gat);
xor XOR2_56 (G236gat, G203gat, G168gat);
xor XOR2_57 (G239gat, G203gat, G171gat);
nand NAND2_58 (G242gat, G1gat, G213gat);
xor XOR2_59 (G243gat, G203gat, G174gat);
nand NAND2_60 (G246gat, G213gat, G11gat);
xor XOR2_61 (G247gat, G203gat, G177gat);
nand NAND2_62 (G250gat, G213gat, G24gat);
xor XOR2_63 (G251gat, G203gat, G180gat);
nand NAND2_64 (G254gat, G213gat, G37gat);
nand NAND2_65 (G255gat, G213gat, G50gat);
nand NAND2_66 (G256gat, G213gat, G63gat);
nand NAND2_67 (G257gat, G213gat, G76gat);
nand NAND2_68 (G258gat, G213gat, G89gat);
nand NAND2_69 (G259gat, G213gat, G102gat);
nand NAND2_70 (G260gat, G224gat, G157gat);
nand NAND2_71 (G263gat, G224gat, G158gat);
nand NAND2_72 (G264gat, G227gat, G183gat);
nand NAND2_73 (G267gat, G230gat, G185gat);
nand NAND2_74 (G270gat, G233gat, G187gat);
nand NAND2_75 (G273gat, G236gat, G189gat);
nand NAND2_76 (G276gat, G239gat, G191gat);
nand NAND2_77 (G279gat, G243gat, G193gat);
nand NAND2_78 (G282gat, G247gat, G195gat);
nand NAND2_79 (G285gat, G251gat, G197gat);
nand NAND2_80 (G288gat, G227gat, G184gat);
nand NAND2_81 (G289gat, G230gat, G186gat);
nand NAND2_82 (G290gat, G233gat, G188gat);
nand NAND2_83 (G291gat, G236gat, G190gat);
nand NAND2_84 (G292gat, G239gat, G192gat);
nand NAND2_85 (G293gat, G243gat, G194gat);
nand NAND2_86 (G294gat, G247gat, G196gat);
nand NAND2_87 (G295gat, G251gat, G198gat);
and AND4_88 (G2950gat, G260gat, G264gat, G267gat, G270gat);
and AND5_89 (G2951gat, G273gat, G276gat, G279gat, G282gat, G285gat);
and AND2_90 (G296gat, G2950gat, G2951gat);
not NOT1_91 (G300gat, G263gat);
not NOT1_92 (G301gat, G288gat);
not NOT1_93 (G302gat, G289gat);
not NOT1_94 (G303gat, G290gat);
not NOT1_95 (G304gat, G291gat);
not NOT1_96 (G305gat, G292gat);
not NOT1_97 (G306gat, G293gat);
not NOT1_98 (G307gat, G294gat);
not NOT1_99 (G308gat, G295gat);
not NOT1_100 (G309gat, G296gat);
not NOT1_101 (G319gat, G296gat);
not NOT1_102 (G329gat, G296gat);
xor XOR2_103 (G330gat, G309gat, G260gat);
xor XOR2_104 (G331gat, G309gat, G264gat);
xor XOR2_105 (G332gat, G309gat, G267gat);
xor XOR2_106 (G333gat, G309gat, G270gat);
nand NAND2_107 (G334gat, G8gat, G319gat);
xor XOR2_108 (G335gat, G309gat, G273gat);
nand NAND2_109 (G336gat, G319gat, G21gat);
xor XOR2_110 (G337gat, G309gat, G276gat);
nand NAND2_111 (G338gat, G319gat, G34gat);
xor XOR2_112 (G339gat, G309gat, G279gat);
nand NAND2_113 (G340gat, G319gat, G47gat);
xor XOR2_114 (G341gat, G309gat, G282gat);
nand NAND2_115 (G342gat, G319gat, G60gat);
xor XOR2_116 (G343gat, G309gat, G285gat);
nand NAND2_117 (G344gat, G319gat, G73gat);
nand NAND2_118 (G345gat, G319gat, G86gat);
nand NAND2_119 (G346gat, G319gat, G99gat);
nand NAND2_120 (G347gat, G319gat, G112gat);
nand NAND2_121 (G348gat, G330gat, G300gat);
nand NAND2_122 (G349gat, G331gat, G301gat);
nand NAND2_123 (G350gat, G332gat, G302gat);
nand NAND2_124 (G351gat, G333gat, G303gat);
nand NAND2_125 (G352gat, G335gat, G304gat);
nand NAND2_126 (G353gat, G337gat, G305gat);
nand NAND2_127 (G354gat, G339gat, G306gat);
nand NAND2_128 (G355gat, G341gat, G307gat);
nand NAND2_129 (G356gat, G343gat, G308gat);
and AND4_130 (G3560gat, G348gat, G349gat, G350gat, G351gat);
and AND5_131 (G3561gat, G352gat, G353gat, G354gat, G355gat, G356gat);
and AND2_132 (G357gat, G3560gat, G3561gat);
not NOT1_133 (G360gat, G357gat);
not NOT1_134 (G370gat, G357gat);
nand NAND2_135 (G371gat, G14gat, G360gat);
nand NAND2_136 (G372gat, G360gat, G27gat);
nand NAND2_137 (G373gat, G360gat, G40gat);
nand NAND2_138 (G374gat, G360gat, G53gat);
nand NAND2_139 (G375gat, G360gat, G66gat);
nand NAND2_140 (G376gat, G360gat, G79gat);
nand NAND2_141 (G377gat, G360gat, G92gat);
nand NAND2_142 (G378gat, G360gat, G105gat);
nand NAND2_143 (G379gat, G360gat, G115gat);
nand NAND4_144 (G380gat, G4gat, G242gat, G334gat, G371gat);
nand NAND4_145 (G381gat, G246gat, G336gat, G372gat, G17gat);
nand NAND4_146 (G386gat, G250gat, G338gat, G373gat, G30gat);
nand NAND4_147 (G393gat, G254gat, G340gat, G374gat, G43gat);
nand NAND4_148 (G399gat, G255gat, G342gat, G375gat, G56gat);
nand NAND4_149 (G404gat, G256gat, G344gat, G376gat, G69gat);
nand NAND4_150 (G407gat, G257gat, G345gat, G377gat, G82gat);
nand NAND4_151 (G411gat, G258gat, G346gat, G378gat, G95gat);
nand NAND4_152 (G414gat, G259gat, G347gat, G379gat, G108gat);
not NOT1_153 (G415gat, G380gat);
and AND4_154 (G4150gat, G381gat, G386gat, G393gat, G399gat);
and AND4_155 (G4151gat, G404gat, G407gat, G411gat, G414gat);
and AND2_156 (G416gat, G4150gat, G4151gat);
not NOT1_157 (G417gat, G393gat);
not NOT1_158 (G418gat, G404gat);
not NOT1_159 (G419gat, G407gat);
not NOT1_160 (G420gat, G411gat);
nor NOR2_161 (G421gat, G415gat, G416gat);
nand NAND2_162 (G422gat, G386gat, G417gat);
nand NAND4_163 (G425gat, G386gat, G393gat, G418gat, G399gat);
nand NAND3_164 (G428gat, G399gat, G393gat, G419gat);
nand NAND4_165 (G429gat, G386gat, G393gat, G407gat, G420gat);
nand NAND4_166 (G430gat, G381gat, G386gat, G422gat, G399gat);
nand NAND4_167 (G431gat, G381gat, G386gat, G425gat, G428gat);
nand NAND4_168 (G432gat, G381gat, G422gat, G425gat, G429gat);

endmodule