module DFF(Q, clk, D);
input D;
input clk;
output Q;
always @(clk)
begin
  Q <= D;
end
endmodule


module c432_libar_24k(G1gat,G4gat,G8gat,G11gat,G14gat,G17gat,G21gat,G24gat,G27gat,G30gat,G34gat,G37gat,G40gat,G43gat,G47gat,G50gat,G53gat,G56gat,G60gat,G63gat,G66gat,G69gat,G73gat,G76gat,G79gat,G82gat,G86gat,G89gat,G92gat,G95gat,G99gat,G102gat,G105gat,G108gat,G112gat,G115gat,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,G223gat,G329gat,G370gat,G421gat,G430gat,G431gat,G432gat);

input G1gat,G4gat,G8gat,G11gat,G14gat,G17gat,G21gat,G24gat,G27gat,G30gat,G34gat,G37gat,G40gat,G43gat,G47gat,G50gat,G53gat,G56gat,G60gat,G63gat,G66gat,G69gat,G73gat,G76gat,G79gat,G82gat,G86gat,G89gat,G92gat,G95gat,G99gat,G102gat,G105gat,G108gat,G112gat,G115gat,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23;
output G223gat,G329gat,G370gat,G421gat,G430gat,G431gat,G432gat;
wire G118gat_enc,G118gat,G119gat_enc,CLK8,LIBAR8,G119gat,G122gat,G123gat_enc,CLK7,LIBAR7,G123gat,G126gat_enc,G126gat,G127gat,G130gat_enc,CLK6,LIBAR6,G130gat,G131gat_enc,G131gat,G134gat,G135gat_enc,CLK5,LIBAR5,G135gat,G138gat_enc,CLK4,LIBAR4,G138gat,G139gat_enc,CLK3,LIBAR3,G139gat,G142gat,G143gat,G146gat,G147gat_enc,CLK2,LIBAR2,G147gat,G150gat_enc,CLK1,LIBAR1,G150gat,G151gat_enc,G151gat,G154gat_enc,G154gat,G157gat_enc,G157gat,G158gat_enc,G158gat,G159gat_enc,G159gat,G162gat_enc,G162gat,G165gat_enc,G165gat,G168gat_enc,G168gat,G171gat,G174gat,G177gat,G180gat,G183gat,G184gat,G185gat_enc,G185gat,G186gat,G187gat_enc,G187gat,G188gat_enc,G188gat,G189gat_enc,G189gat,G190gat_enc,G190gat,G191gat,G192gat,G193gat,G194gat,G195gat,G196gat,G197gat,G198gat,G1980gat,G1981gat,G199gat,G203gat,G213gat,G224gat,G227gat,G230gat,G233gat,G236gat,G239gat,G242gat,G243gat,G246gat,G247gat,G250gat,G251gat,G254gat,G255gat,G256gat,G257gat,G258gat,G259gat,G260gat,G263gat,G264gat,G267gat,G270gat,G273gat,G276gat,G279gat,G282gat,G285gat,G288gat,G289gat,G290gat,G291gat,G292gat,G293gat,G294gat,G295gat,G2950gat,G2951gat,G296gat,G300gat,G301gat,G302gat,G303gat,G304gat,G305gat,G306gat,G307gat,G308gat,G309gat,G319gat,G330gat,G331gat,G332gat,G333gat,G334gat,G335gat,G336gat,G337gat,G338gat,G339gat,G340gat,G341gat,G342gat,G343gat,G344gat,G345gat,G346gat,G347gat,G348gat,G349gat,G350gat,G351gat,G352gat,G353gat,G354gat,G355gat,G356gat,G3560gat,G3561gat,G357gat,G360gat,G371gat,G372gat,G373gat,G374gat,G375gat,G376gat,G377gat,G378gat,G379gat,G380gat,G381gat,G386gat,G393gat,G399gat,G404gat,G407gat,G411gat,G414gat,G415gat,G4150gat,G4151gat,G416gat,G417gat,G418gat,G419gat,G420gat,G422gat,G425gat,G428gat,G429gat;

not NOT1_1 (G118gat_enc, G1gat);
xor XOR2_2 (G118gat, keyinput0, G118gat_enc);
not NOT1_3 (G119gat_enc, G4gat);
nor NOR2_4 (CLK8, G119gat_enc, G118gat);
dff DFF2_5 (LIBAR8, CLK8, keyinput1);
xor XOR2_6 (G119gat, LIBAR8, G119gat_enc);
not NOT1_7 (G122gat, G11gat);
not NOT1_8 (G123gat_enc, G17gat);
nor NOR2_9 (CLK7, G123gat_enc, G122gat);
dff DFF2_10 (LIBAR7, CLK7, keyinput2);
xnor XNOR2_11 (G123gat, LIBAR7, G123gat_enc);
not NOT1_12 (G126gat_enc, G24gat);
xor XOR2_13 (G126gat, keyinput3, G126gat_enc);
not NOT1_14 (G127gat, G30gat);
not NOT1_15 (G130gat_enc, G37gat);
nor NOR2_16 (CLK6, G130gat_enc, G127gat);
dff DFF2_17 (LIBAR6, CLK6, keyinput4);
xnor XNOR2_18 (G130gat, LIBAR6, G130gat_enc);
not NOT1_19 (G131gat_enc, G43gat);
xor XOR2_20 (G131gat, keyinput5, G131gat_enc);
not NOT1_21 (G134gat, G50gat);
not NOT1_22 (G135gat_enc, G56gat);
nor NOR2_23 (CLK5, G135gat_enc, G134gat);
dff DFF2_24 (LIBAR5, CLK5, keyinput6);
xnor XNOR2_25 (G135gat, LIBAR5, G135gat_enc);
not NOT1_26 (G138gat_enc, G63gat);
nor NOR2_27 (CLK4, G138gat_enc, G135gat);
dff DFF2_28 (LIBAR4, CLK4, keyinput7);
xor XOR2_29 (G138gat, LIBAR4, G138gat_enc);
not NOT1_30 (G139gat_enc, G69gat);
nor NOR2_31 (CLK3, G139gat_enc, G138gat);
dff DFF2_32 (LIBAR3, CLK3, keyinput8);
xnor XNOR2_33 (G139gat, LIBAR3, G139gat_enc);
not NOT1_34 (G142gat, G76gat);
not NOT1_35 (G143gat, G82gat);
not NOT1_36 (G146gat, G89gat);
not NOT1_37 (G147gat_enc, G95gat);
nor NOR2_38 (CLK2, G147gat_enc, G146gat);
dff DFF2_39 (LIBAR2, CLK2, keyinput9);
xnor XNOR2_40 (G147gat, LIBAR2, G147gat_enc);
not NOT1_41 (G150gat_enc, G102gat);
nor NOR2_42 (CLK1, G150gat_enc, G147gat);
dff DFF2_43 (LIBAR1, CLK1, keyinput10);
xnor XNOR2_44 (G150gat, LIBAR1, G150gat_enc);
not NOT1_45 (G151gat_enc, G108gat);
xnor XNOR2_46 (G151gat, keyinput11, G151gat_enc);
nand NAND2_47 (G154gat_enc, G118gat, G4gat);
xor XOR2_48 (G154gat, keyinput12, G154gat_enc);
nor NOR2_49 (G157gat_enc, G8gat, G119gat);
xor XOR2_50 (G157gat, keyinput13, G157gat_enc);
nor NOR2_51 (G158gat_enc, G14gat, G119gat);
xor XOR2_52 (G158gat, keyinput14, G158gat_enc);
nand NAND2_53 (G159gat_enc, G122gat, G17gat);
xnor XNOR2_54 (G159gat, keyinput15, G159gat_enc);
nand NAND2_55 (G162gat_enc, G126gat, G30gat);
xor XOR2_56 (G162gat, keyinput16, G162gat_enc);
nand NAND2_57 (G165gat_enc, G130gat, G43gat);
xnor XNOR2_58 (G165gat, keyinput17, G165gat_enc);
nand NAND2_59 (G168gat_enc, G134gat, G56gat);
xor XOR2_60 (G168gat, keyinput18, G168gat_enc);
nand NAND2_61 (G171gat, G138gat, G69gat);
nand NAND2_62 (G174gat, G142gat, G82gat);
nand NAND2_63 (G177gat, G146gat, G95gat);
nand NAND2_64 (G180gat, G150gat, G108gat);
nor NOR2_65 (G183gat, G21gat, G123gat);
nor NOR2_66 (G184gat, G27gat, G123gat);
nor NOR2_67 (G185gat_enc, G34gat, G127gat);
xnor XNOR2_68 (G185gat, keyinput19, G185gat_enc);
nor NOR2_69 (G186gat, G40gat, G127gat);
nor NOR2_70 (G187gat_enc, G47gat, G131gat);
xnor XNOR2_71 (G187gat, keyinput20, G187gat_enc);
nor NOR2_72 (G188gat_enc, G53gat, G131gat);
xnor XNOR2_73 (G188gat, keyinput21, G188gat_enc);
nor NOR2_74 (G189gat_enc, G60gat, G135gat);
xor XOR2_75 (G189gat, keyinput22, G189gat_enc);
nor NOR2_76 (G190gat_enc, G66gat, G135gat);
xnor XNOR2_77 (G190gat, keyinput23, G190gat_enc);
nor NOR2_78 (G191gat, G73gat, G139gat);
nor NOR2_79 (G192gat, G79gat, G139gat);
nor NOR2_80 (G193gat, G86gat, G143gat);
nor NOR2_81 (G194gat, G92gat, G143gat);
nor NOR2_82 (G195gat, G99gat, G147gat);
nor NOR2_83 (G196gat, G105gat, G147gat);
nor NOR2_84 (G197gat, G112gat, G151gat);
nor NOR2_85 (G198gat, G115gat, G151gat);
and AND4_86 (G1980gat, G154gat, G159gat, G162gat, G165gat);
and AND5_87 (G1981gat, G168gat, G171gat, G174gat, G177gat, G180gat);
and AND2_88 (G199gat, G1980gat, G1981gat);
not NOT1_89 (G203gat, G199gat);
not NOT1_90 (G213gat, G199gat);
not NOT1_91 (G223gat, G199gat);
xor XOR2_92 (G224gat, G203gat, G154gat);
xor XOR2_93 (G227gat, G203gat, G159gat);
xor XOR2_94 (G230gat, G203gat, G162gat);
xor XOR2_95 (G233gat, G203gat, G165gat);
xor XOR2_96 (G236gat, G203gat, G168gat);
xor XOR2_97 (G239gat, G203gat, G171gat);
nand NAND2_98 (G242gat, G1gat, G213gat);
xor XOR2_99 (G243gat, G203gat, G174gat);
nand NAND2_100 (G246gat, G213gat, G11gat);
xor XOR2_101 (G247gat, G203gat, G177gat);
nand NAND2_102 (G250gat, G213gat, G24gat);
xor XOR2_103 (G251gat, G203gat, G180gat);
nand NAND2_104 (G254gat, G213gat, G37gat);
nand NAND2_105 (G255gat, G213gat, G50gat);
nand NAND2_106 (G256gat, G213gat, G63gat);
nand NAND2_107 (G257gat, G213gat, G76gat);
nand NAND2_108 (G258gat, G213gat, G89gat);
nand NAND2_109 (G259gat, G213gat, G102gat);
nand NAND2_110 (G260gat, G224gat, G157gat);
nand NAND2_111 (G263gat, G224gat, G158gat);
nand NAND2_112 (G264gat, G227gat, G183gat);
nand NAND2_113 (G267gat, G230gat, G185gat);
nand NAND2_114 (G270gat, G233gat, G187gat);
nand NAND2_115 (G273gat, G236gat, G189gat);
nand NAND2_116 (G276gat, G239gat, G191gat);
nand NAND2_117 (G279gat, G243gat, G193gat);
nand NAND2_118 (G282gat, G247gat, G195gat);
nand NAND2_119 (G285gat, G251gat, G197gat);
nand NAND2_120 (G288gat, G227gat, G184gat);
nand NAND2_121 (G289gat, G230gat, G186gat);
nand NAND2_122 (G290gat, G233gat, G188gat);
nand NAND2_123 (G291gat, G236gat, G190gat);
nand NAND2_124 (G292gat, G239gat, G192gat);
nand NAND2_125 (G293gat, G243gat, G194gat);
nand NAND2_126 (G294gat, G247gat, G196gat);
nand NAND2_127 (G295gat, G251gat, G198gat);
and AND4_128 (G2950gat, G260gat, G264gat, G267gat, G270gat);
and AND5_129 (G2951gat, G273gat, G276gat, G279gat, G282gat, G285gat);
and AND2_130 (G296gat, G2950gat, G2951gat);
not NOT1_131 (G300gat, G263gat);
not NOT1_132 (G301gat, G288gat);
not NOT1_133 (G302gat, G289gat);
not NOT1_134 (G303gat, G290gat);
not NOT1_135 (G304gat, G291gat);
not NOT1_136 (G305gat, G292gat);
not NOT1_137 (G306gat, G293gat);
not NOT1_138 (G307gat, G294gat);
not NOT1_139 (G308gat, G295gat);
not NOT1_140 (G309gat, G296gat);
not NOT1_141 (G319gat, G296gat);
not NOT1_142 (G329gat, G296gat);
xor XOR2_143 (G330gat, G309gat, G260gat);
xor XOR2_144 (G331gat, G309gat, G264gat);
xor XOR2_145 (G332gat, G309gat, G267gat);
xor XOR2_146 (G333gat, G309gat, G270gat);
nand NAND2_147 (G334gat, G8gat, G319gat);
xor XOR2_148 (G335gat, G309gat, G273gat);
nand NAND2_149 (G336gat, G319gat, G21gat);
xor XOR2_150 (G337gat, G309gat, G276gat);
nand NAND2_151 (G338gat, G319gat, G34gat);
xor XOR2_152 (G339gat, G309gat, G279gat);
nand NAND2_153 (G340gat, G319gat, G47gat);
xor XOR2_154 (G341gat, G309gat, G282gat);
nand NAND2_155 (G342gat, G319gat, G60gat);
xor XOR2_156 (G343gat, G309gat, G285gat);
nand NAND2_157 (G344gat, G319gat, G73gat);
nand NAND2_158 (G345gat, G319gat, G86gat);
nand NAND2_159 (G346gat, G319gat, G99gat);
nand NAND2_160 (G347gat, G319gat, G112gat);
nand NAND2_161 (G348gat, G330gat, G300gat);
nand NAND2_162 (G349gat, G331gat, G301gat);
nand NAND2_163 (G350gat, G332gat, G302gat);
nand NAND2_164 (G351gat, G333gat, G303gat);
nand NAND2_165 (G352gat, G335gat, G304gat);
nand NAND2_166 (G353gat, G337gat, G305gat);
nand NAND2_167 (G354gat, G339gat, G306gat);
nand NAND2_168 (G355gat, G341gat, G307gat);
nand NAND2_169 (G356gat, G343gat, G308gat);
and AND4_170 (G3560gat, G348gat, G349gat, G350gat, G351gat);
and AND5_171 (G3561gat, G352gat, G353gat, G354gat, G355gat, G356gat);
and AND2_172 (G357gat, G3560gat, G3561gat);
not NOT1_173 (G360gat, G357gat);
not NOT1_174 (G370gat, G357gat);
nand NAND2_175 (G371gat, G14gat, G360gat);
nand NAND2_176 (G372gat, G360gat, G27gat);
nand NAND2_177 (G373gat, G360gat, G40gat);
nand NAND2_178 (G374gat, G360gat, G53gat);
nand NAND2_179 (G375gat, G360gat, G66gat);
nand NAND2_180 (G376gat, G360gat, G79gat);
nand NAND2_181 (G377gat, G360gat, G92gat);
nand NAND2_182 (G378gat, G360gat, G105gat);
nand NAND2_183 (G379gat, G360gat, G115gat);
nand NAND4_184 (G380gat, G4gat, G242gat, G334gat, G371gat);
nand NAND4_185 (G381gat, G246gat, G336gat, G372gat, G17gat);
nand NAND4_186 (G386gat, G250gat, G338gat, G373gat, G30gat);
nand NAND4_187 (G393gat, G254gat, G340gat, G374gat, G43gat);
nand NAND4_188 (G399gat, G255gat, G342gat, G375gat, G56gat);
nand NAND4_189 (G404gat, G256gat, G344gat, G376gat, G69gat);
nand NAND4_190 (G407gat, G257gat, G345gat, G377gat, G82gat);
nand NAND4_191 (G411gat, G258gat, G346gat, G378gat, G95gat);
nand NAND4_192 (G414gat, G259gat, G347gat, G379gat, G108gat);
not NOT1_193 (G415gat, G380gat);
and AND4_194 (G4150gat, G381gat, G386gat, G393gat, G399gat);
and AND4_195 (G4151gat, G404gat, G407gat, G411gat, G414gat);
and AND2_196 (G416gat, G4150gat, G4151gat);
not NOT1_197 (G417gat, G393gat);
not NOT1_198 (G418gat, G404gat);
not NOT1_199 (G419gat, G407gat);
not NOT1_200 (G420gat, G411gat);
nor NOR2_201 (G421gat, G415gat, G416gat);
nand NAND2_202 (G422gat, G386gat, G417gat);
nand NAND4_203 (G425gat, G386gat, G393gat, G418gat, G399gat);
nand NAND3_204 (G428gat, G399gat, G393gat, G419gat);
nand NAND4_205 (G429gat, G386gat, G393gat, G407gat, G420gat);
nand NAND4_206 (G430gat, G381gat, G386gat, G422gat, G399gat);
nand NAND4_207 (G431gat, G381gat, G386gat, G425gat, G428gat);
nand NAND4_208 (G432gat, G381gat, G422gat, G425gat, G429gat);

endmodule