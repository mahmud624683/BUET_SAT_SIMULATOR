module c432_rll_32k(G1gat,G4gat,G8gat,G11gat,G14gat,G17gat,G21gat,G24gat,G27gat,G30gat,G34gat,G37gat,G40gat,G43gat,G47gat,G50gat,G53gat,G56gat,G60gat,G63gat,G66gat,G69gat,G73gat,G76gat,G79gat,G82gat,G86gat,G89gat,G92gat,G95gat,G99gat,G102gat,G105gat,G108gat,G112gat,G115gat,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,G223gat,G329gat,G370gat,G421gat,G430gat,G431gat,G432gat);

input G1gat,G4gat,G8gat,G11gat,G14gat,G17gat,G21gat,G24gat,G27gat,G30gat,G34gat,G37gat,G40gat,G43gat,G47gat,G50gat,G53gat,G56gat,G60gat,G63gat,G66gat,G69gat,G73gat,G76gat,G79gat,G82gat,G86gat,G89gat,G92gat,G95gat,G99gat,G102gat,G105gat,G108gat,G112gat,G115gat,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31;
output G223gat,G329gat,G370gat,G421gat,G430gat,G431gat,G432gat;
wire G118gat,G119gat_enc,G119gat,G122gat_enc,G122gat,G123gat_enc,G123gat,G126gat,G127gat_enc,G127gat,G130gat,G131gat_enc,G131gat,G134gat_enc,G134gat,G135gat_enc,G135gat,G138gat_enc,G138gat,G139gat_enc,G139gat,G142gat,G143gat_enc,G143gat,G146gat_enc,G146gat,G147gat,G150gat_enc,G150gat,G151gat,G154gat,G157gat,G158gat,G159gat,G162gat_enc,G162gat,G165gat_enc,G165gat,G168gat,G171gat_enc,G171gat,G174gat_enc,G174gat,G177gat,G180gat,G183gat_enc,G183gat,G184gat_enc,G184gat,G185gat_enc,G185gat,G186gat_enc,G186gat,G187gat,G188gat,G189gat_enc,G189gat,G190gat,G191gat,G192gat,G193gat_enc,G193gat,G194gat_enc,G194gat,G195gat,G196gat,G197gat_enc,G197gat,G198gat_enc,G198gat,G1980gat,G1981gat_enc,G1981gat,G199gat_enc,G199gat,G203gat_enc,G203gat,G213gat_enc,G213gat,G224gat,G227gat_enc,G227gat,G230gat_enc,G230gat,G233gat,G236gat,G239gat,G242gat,G243gat,G246gat,G247gat,G250gat,G251gat,G254gat_enc,G254gat,G255gat,G256gat,G257gat,G258gat,G259gat,G260gat,G263gat,G264gat,G267gat,G270gat,G273gat,G276gat,G279gat,G282gat,G285gat,G288gat,G289gat,G290gat,G291gat,G292gat,G293gat,G294gat,G295gat,G2950gat,G2951gat,G296gat,G300gat,G301gat,G302gat,G303gat,G304gat,G305gat,G306gat,G307gat,G308gat,G309gat,G319gat,G330gat,G331gat,G332gat,G333gat,G334gat,G335gat,G336gat,G337gat,G338gat,G339gat,G340gat,G341gat,G342gat,G343gat,G344gat,G345gat,G346gat,G347gat,G348gat,G349gat,G350gat,G351gat,G352gat,G353gat,G354gat,G355gat,G356gat,G3560gat,G3561gat,G357gat,G360gat,G371gat,G372gat,G373gat,G374gat,G375gat,G376gat,G377gat,G378gat,G379gat,G380gat,G381gat,G386gat,G393gat,G399gat,G404gat,G407gat,G411gat,G414gat,G415gat,G4150gat,G4151gat,G416gat,G417gat,G418gat,G419gat,G420gat,G422gat,G425gat,G428gat,G429gat;

not NOT1_1 (G118gat, G1gat);
not NOT1_2 (G119gat_enc, G4gat);
xnor XNOR2_3 (G119gat, keyinput0, G119gat_enc);
not NOT1_4 (G122gat_enc, G11gat);
xor XOR2_5 (G122gat, keyinput1, G122gat_enc);
not NOT1_6 (G123gat_enc, G17gat);
xor XOR2_7 (G123gat, keyinput2, G123gat_enc);
not NOT1_8 (G126gat, G24gat);
not NOT1_9 (G127gat_enc, G30gat);
xnor XNOR2_10 (G127gat, keyinput3, G127gat_enc);
not NOT1_11 (G130gat, G37gat);
not NOT1_12 (G131gat_enc, G43gat);
xnor XNOR2_13 (G131gat, keyinput4, G131gat_enc);
not NOT1_14 (G134gat_enc, G50gat);
xor XOR2_15 (G134gat, keyinput5, G134gat_enc);
not NOT1_16 (G135gat_enc, G56gat);
xor XOR2_17 (G135gat, keyinput6, G135gat_enc);
not NOT1_18 (G138gat_enc, G63gat);
xor XOR2_19 (G138gat, keyinput7, G138gat_enc);
not NOT1_20 (G139gat_enc, G69gat);
xnor XNOR2_21 (G139gat, keyinput8, G139gat_enc);
not NOT1_22 (G142gat, G76gat);
not NOT1_23 (G143gat_enc, G82gat);
xnor XNOR2_24 (G143gat, keyinput9, G143gat_enc);
not NOT1_25 (G146gat_enc, G89gat);
xnor XNOR2_26 (G146gat, keyinput10, G146gat_enc);
not NOT1_27 (G147gat, G95gat);
not NOT1_28 (G150gat_enc, G102gat);
xnor XNOR2_29 (G150gat, keyinput11, G150gat_enc);
not NOT1_30 (G151gat, G108gat);
nand NAND2_31 (G154gat, G118gat, G4gat);
nor NOR2_32 (G157gat, G8gat, G119gat);
nor NOR2_33 (G158gat, G14gat, G119gat);
nand NAND2_34 (G159gat, G122gat, G17gat);
nand NAND2_35 (G162gat_enc, G126gat, G30gat);
xnor XNOR2_36 (G162gat, keyinput12, G162gat_enc);
nand NAND2_37 (G165gat_enc, G130gat, G43gat);
xor XOR2_38 (G165gat, keyinput13, G165gat_enc);
nand NAND2_39 (G168gat, G134gat, G56gat);
nand NAND2_40 (G171gat_enc, G138gat, G69gat);
xnor XNOR2_41 (G171gat, keyinput14, G171gat_enc);
nand NAND2_42 (G174gat_enc, G142gat, G82gat);
xor XOR2_43 (G174gat, keyinput15, G174gat_enc);
nand NAND2_44 (G177gat, G146gat, G95gat);
nand NAND2_45 (G180gat, G150gat, G108gat);
nor NOR2_46 (G183gat_enc, G21gat, G123gat);
xnor XNOR2_47 (G183gat, keyinput16, G183gat_enc);
nor NOR2_48 (G184gat_enc, G27gat, G123gat);
xor XOR2_49 (G184gat, keyinput17, G184gat_enc);
nor NOR2_50 (G185gat_enc, G34gat, G127gat);
xnor XNOR2_51 (G185gat, keyinput18, G185gat_enc);
nor NOR2_52 (G186gat_enc, G40gat, G127gat);
xor XOR2_53 (G186gat, keyinput19, G186gat_enc);
nor NOR2_54 (G187gat, G47gat, G131gat);
nor NOR2_55 (G188gat, G53gat, G131gat);
nor NOR2_56 (G189gat_enc, G60gat, G135gat);
xnor XNOR2_57 (G189gat, keyinput20, G189gat_enc);
nor NOR2_58 (G190gat, G66gat, G135gat);
nor NOR2_59 (G191gat, G73gat, G139gat);
nor NOR2_60 (G192gat, G79gat, G139gat);
nor NOR2_61 (G193gat_enc, G86gat, G143gat);
xnor XNOR2_62 (G193gat, keyinput21, G193gat_enc);
nor NOR2_63 (G194gat_enc, G92gat, G143gat);
xnor XNOR2_64 (G194gat, keyinput22, G194gat_enc);
nor NOR2_65 (G195gat, G99gat, G147gat);
nor NOR2_66 (G196gat, G105gat, G147gat);
nor NOR2_67 (G197gat_enc, G112gat, G151gat);
xnor XNOR2_68 (G197gat, keyinput23, G197gat_enc);
nor NOR2_69 (G198gat_enc, G115gat, G151gat);
xor XOR2_70 (G198gat, keyinput24, G198gat_enc);
and AND4_71 (G1980gat, G154gat, G159gat, G162gat, G165gat);
and AND5_72 (G1981gat_enc, G168gat, G171gat, G174gat, G177gat, G180gat);
xnor XNOR2_73 (G1981gat, keyinput25, G1981gat_enc);
and AND2_74 (G199gat_enc, G1980gat, G1981gat);
xor XOR2_75 (G199gat, keyinput26, G199gat_enc);
not NOT1_76 (G203gat_enc, G199gat);
xnor XNOR2_77 (G203gat, keyinput27, G203gat_enc);
not NOT1_78 (G213gat_enc, G199gat);
xor XOR2_79 (G213gat, keyinput28, G213gat_enc);
not NOT1_80 (G223gat, G199gat);
xor XOR2_81 (G224gat, G203gat, G154gat);
xor XOR2_82 (G227gat_enc, G203gat, G159gat);
xnor XNOR2_83 (G227gat, keyinput29, G227gat_enc);
xor XOR2_84 (G230gat_enc, G203gat, G162gat);
xor XOR2_85 (G230gat, keyinput30, G230gat_enc);
xor XOR2_86 (G233gat, G203gat, G165gat);
xor XOR2_87 (G236gat, G203gat, G168gat);
xor XOR2_88 (G239gat, G203gat, G171gat);
nand NAND2_89 (G242gat, G1gat, G213gat);
xor XOR2_90 (G243gat, G203gat, G174gat);
nand NAND2_91 (G246gat, G213gat, G11gat);
xor XOR2_92 (G247gat, G203gat, G177gat);
nand NAND2_93 (G250gat, G213gat, G24gat);
xor XOR2_94 (G251gat, G203gat, G180gat);
nand NAND2_95 (G254gat_enc, G213gat, G37gat);
xnor XNOR2_96 (G254gat, keyinput31, G254gat_enc);
nand NAND2_97 (G255gat, G213gat, G50gat);
nand NAND2_98 (G256gat, G213gat, G63gat);
nand NAND2_99 (G257gat, G213gat, G76gat);
nand NAND2_100 (G258gat, G213gat, G89gat);
nand NAND2_101 (G259gat, G213gat, G102gat);
nand NAND2_102 (G260gat, G224gat, G157gat);
nand NAND2_103 (G263gat, G224gat, G158gat);
nand NAND2_104 (G264gat, G227gat, G183gat);
nand NAND2_105 (G267gat, G230gat, G185gat);
nand NAND2_106 (G270gat, G233gat, G187gat);
nand NAND2_107 (G273gat, G236gat, G189gat);
nand NAND2_108 (G276gat, G239gat, G191gat);
nand NAND2_109 (G279gat, G243gat, G193gat);
nand NAND2_110 (G282gat, G247gat, G195gat);
nand NAND2_111 (G285gat, G251gat, G197gat);
nand NAND2_112 (G288gat, G227gat, G184gat);
nand NAND2_113 (G289gat, G230gat, G186gat);
nand NAND2_114 (G290gat, G233gat, G188gat);
nand NAND2_115 (G291gat, G236gat, G190gat);
nand NAND2_116 (G292gat, G239gat, G192gat);
nand NAND2_117 (G293gat, G243gat, G194gat);
nand NAND2_118 (G294gat, G247gat, G196gat);
nand NAND2_119 (G295gat, G251gat, G198gat);
and AND4_120 (G2950gat, G260gat, G264gat, G267gat, G270gat);
and AND5_121 (G2951gat, G273gat, G276gat, G279gat, G282gat, G285gat);
and AND2_122 (G296gat, G2950gat, G2951gat);
not NOT1_123 (G300gat, G263gat);
not NOT1_124 (G301gat, G288gat);
not NOT1_125 (G302gat, G289gat);
not NOT1_126 (G303gat, G290gat);
not NOT1_127 (G304gat, G291gat);
not NOT1_128 (G305gat, G292gat);
not NOT1_129 (G306gat, G293gat);
not NOT1_130 (G307gat, G294gat);
not NOT1_131 (G308gat, G295gat);
not NOT1_132 (G309gat, G296gat);
not NOT1_133 (G319gat, G296gat);
not NOT1_134 (G329gat, G296gat);
xor XOR2_135 (G330gat, G309gat, G260gat);
xor XOR2_136 (G331gat, G309gat, G264gat);
xor XOR2_137 (G332gat, G309gat, G267gat);
xor XOR2_138 (G333gat, G309gat, G270gat);
nand NAND2_139 (G334gat, G8gat, G319gat);
xor XOR2_140 (G335gat, G309gat, G273gat);
nand NAND2_141 (G336gat, G319gat, G21gat);
xor XOR2_142 (G337gat, G309gat, G276gat);
nand NAND2_143 (G338gat, G319gat, G34gat);
xor XOR2_144 (G339gat, G309gat, G279gat);
nand NAND2_145 (G340gat, G319gat, G47gat);
xor XOR2_146 (G341gat, G309gat, G282gat);
nand NAND2_147 (G342gat, G319gat, G60gat);
xor XOR2_148 (G343gat, G309gat, G285gat);
nand NAND2_149 (G344gat, G319gat, G73gat);
nand NAND2_150 (G345gat, G319gat, G86gat);
nand NAND2_151 (G346gat, G319gat, G99gat);
nand NAND2_152 (G347gat, G319gat, G112gat);
nand NAND2_153 (G348gat, G330gat, G300gat);
nand NAND2_154 (G349gat, G331gat, G301gat);
nand NAND2_155 (G350gat, G332gat, G302gat);
nand NAND2_156 (G351gat, G333gat, G303gat);
nand NAND2_157 (G352gat, G335gat, G304gat);
nand NAND2_158 (G353gat, G337gat, G305gat);
nand NAND2_159 (G354gat, G339gat, G306gat);
nand NAND2_160 (G355gat, G341gat, G307gat);
nand NAND2_161 (G356gat, G343gat, G308gat);
and AND4_162 (G3560gat, G348gat, G349gat, G350gat, G351gat);
and AND5_163 (G3561gat, G352gat, G353gat, G354gat, G355gat, G356gat);
and AND2_164 (G357gat, G3560gat, G3561gat);
not NOT1_165 (G360gat, G357gat);
not NOT1_166 (G370gat, G357gat);
nand NAND2_167 (G371gat, G14gat, G360gat);
nand NAND2_168 (G372gat, G360gat, G27gat);
nand NAND2_169 (G373gat, G360gat, G40gat);
nand NAND2_170 (G374gat, G360gat, G53gat);
nand NAND2_171 (G375gat, G360gat, G66gat);
nand NAND2_172 (G376gat, G360gat, G79gat);
nand NAND2_173 (G377gat, G360gat, G92gat);
nand NAND2_174 (G378gat, G360gat, G105gat);
nand NAND2_175 (G379gat, G360gat, G115gat);
nand NAND4_176 (G380gat, G4gat, G242gat, G334gat, G371gat);
nand NAND4_177 (G381gat, G246gat, G336gat, G372gat, G17gat);
nand NAND4_178 (G386gat, G250gat, G338gat, G373gat, G30gat);
nand NAND4_179 (G393gat, G254gat, G340gat, G374gat, G43gat);
nand NAND4_180 (G399gat, G255gat, G342gat, G375gat, G56gat);
nand NAND4_181 (G404gat, G256gat, G344gat, G376gat, G69gat);
nand NAND4_182 (G407gat, G257gat, G345gat, G377gat, G82gat);
nand NAND4_183 (G411gat, G258gat, G346gat, G378gat, G95gat);
nand NAND4_184 (G414gat, G259gat, G347gat, G379gat, G108gat);
not NOT1_185 (G415gat, G380gat);
and AND4_186 (G4150gat, G381gat, G386gat, G393gat, G399gat);
and AND4_187 (G4151gat, G404gat, G407gat, G411gat, G414gat);
and AND2_188 (G416gat, G4150gat, G4151gat);
not NOT1_189 (G417gat, G393gat);
not NOT1_190 (G418gat, G404gat);
not NOT1_191 (G419gat, G407gat);
not NOT1_192 (G420gat, G411gat);
nor NOR2_193 (G421gat, G415gat, G416gat);
nand NAND2_194 (G422gat, G386gat, G417gat);
nand NAND4_195 (G425gat, G386gat, G393gat, G418gat, G399gat);
nand NAND3_196 (G428gat, G399gat, G393gat, G419gat);
nand NAND4_197 (G429gat, G386gat, G393gat, G407gat, G420gat);
nand NAND4_198 (G430gat, G381gat, G386gat, G422gat, G399gat);
nand NAND4_199 (G431gat, G381gat, G386gat, G425gat, G428gat);
nand NAND4_200 (G432gat, G381gat, G422gat, G425gat, G429gat);

endmodule