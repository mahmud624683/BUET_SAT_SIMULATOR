module cac32k(n1,n18,n35,n52,n69,n86,n103,n120,n137,n154,n171,n188,n205,n222,n239,n256,n273,n290,n307,n324,n341,n358,n375,n392,n409,n426,n443,n460,n477,n494,n511,n528,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,n545,n1581,n1901,n2223,n2548,n2877,n3211,n3552,n3895,n4241,n4591,n4946,n5308,n5672,n5971,n6123,n6150,n6160,n6170,n6180,n6190,n6200,n6210,n6220,n6230,n6240,n6250,n6260,n6270,n6280,n6287,n6288);

input n1,n18,n35,n52,n69,n86,n103,n120,n137,n154,n171,n188,n205,n222,n239,n256,n273,n290,n307,n324,n341,n358,n375,n392,n409,n426,n443,n460,n477,n494,n511,n528,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31;
output n545,n1581,n1901,n2223,n2548,n2877,n3211,n3552,n3895,n4241,n4591,n4946,n5308,n5672,n5971,n6123,n6150,n6160,n6170,n6180,n6190,n6200,n6210,n6220,n6230,n6240,n6250,n6260,n6270,n6280,n6287,n6288;
wire wire81,wire163,wire252,wire341,wire428,wire510,wire590,wire691,wire769,wire866,wire949,wire1039,wire1129,wire1315,wire1319,wire1323,wire1325,wire1327,wire1331,wire1335,wire1339,wire1343,wire1347,wire1351,wire1353,wire1355,wire1365,wire1369,wire1371,wire1373,wire1375,wire1377,wire1381,wire1385,wire1389,wire1393,wire1397,wire1409,wire1410,wire1413,wire1414,wire1417,wire1418,wire1421,wire1422,wire1425,wire1426,wire1429,wire1430,wire1500,wire1501,wire1504,wire1505,wire1578,wire1579,wire1580,wire1581,wire1582,wire1583,wire1584,wire1585,wire1586,wire1587,wire1588,wire1589,wire1590,wire1591,wire1592,wire1593,wire1594,wire1595,wire1596,wire1597,wire1598,wire1599,wire1600,wire1601,wire1602,wire1603,wire1604,wire1605,wire1606,wire1607,wire1608,wire1609,wire1610,wire1611,wire1612,wire1613,wire1614,wire1615,wire1616,wire1617,wire1618,wire1619,wire1620,wire1621,wire1622,wire1623,wire1624,wire1625,wire1626,wire1627,wire1628,wire1629,wire1630,wire1631,wire1632,wire1633,wire1634,wire1635,wire1636,wire1637,wire1638,wire1639,wire1640,wire1641,wire1642,wire1643,wire1644,wire1645,wire1646,wire1647,wire1648,wire1649,wire1650,wire1651,wire1652,wire1653,wire1654,wire1655,wire1656,wire1657,wire1658,wire1659,wire1660,wire1661,wire1662,wire1663,wire1664,wire1665,wire1666,wire1667,n_67,n_4,n_5,n_29,n_12,n_13,n_15,n_26,n_21,n_27,n_73,n_19,n_20,n_22,n_31,n_1,n_0,n_8,n_9,n_16,n_23,n_24,n_25,n_28,n_11,n_14,n_30,n_17,n_89,n_18,n_87,n_77,wire1668,wire1669,wire1670,wire1672,wire1673,wire1674,wire1304,wire1305,wire1308,wire1309,wire1316,wire1317,wire1320,wire1321,wire1324,wire1328,wire1329,wire1332,wire1333,wire1336,wire1337,wire1340,wire1341,wire1344,wire1345,wire1348,wire1349,wire1352,wire1356,wire1357,wire1366,wire1367,wire1370,wire1374,wire1378,wire1379,wire1382,wire1383,wire1386,wire1387,wire1390,wire1391,wire1394,wire1395,wire1398,wire1399,wire1411,wire1415,wire1419,wire1423,wire1427,wire1431,wire1433,wire1434,wire1435,wire1436,wire1437,wire1438,wire1439,wire1440,wire1441,wire1442,wire1443,wire1444,wire1445,wire1446,wire1447,wire1448,wire1449,wire1450,wire1451,wire1452,wire1453,wire1454,wire1455,wire1456,wire1457,wire1458,wire1459,wire1460,wire1461,wire1462,wire1463,wire1464,wire1465,wire1466,wire1467,wire1468,wire1469,wire1470,wire1471,wire1472,wire1473,wire1474,wire1475,wire1476,wire1477,wire1478,wire1479,wire1480,wire1481,wire1482,wire1483,wire1484,wire1485,wire1486,wire1487,wire1488,wire1489,wire1490,wire1491,wire1492,wire1493,wire1494,wire1495,wire1496,wire1497,wire1498,wire1499,wire1502,wire1506,wire1508,wire1509,wire1510,wire1511,wire1512,wire1513,wire1514,wire1515,wire1516,wire1517,wire1518,wire1519,wire1520,wire1521,wire1522,wire1523,wire1524,wire1525,wire1526,wire1527,wire1528,wire1529,wire1530,wire1531,wire1532,wire1533,wire1534,wire1535,wire1536,wire1537,wire1538,wire1539,wire1540,wire1541,wire1542,wire1543,wire1544,wire1545,wire1546,wire1547,wire1548,wire1549,wire1550,wire1551,wire1552,wire1553,wire1554,wire1555,wire1556,wire1557,wire1558,wire1559,wire1560,wire1561,wire1562,wire1563,wire1564,wire1565,wire1566,wire1567,wire1568,wire1569,wire1570,wire1571,wire1572,wire1573,wire1574,wire1575,wire1576,wire1577,n_63,n_639,n_47,n_1168,n_1159,n_729,n_58,n_127,n_903,n_255,n_44,n_727,n_868,n_552,n_463,n_1079,n_269,n_567,n_760,n_60,n_956,n_1175,n_962,n_1179,n_161,n_992,n_41,n_919,n_930,n_1245,n_1448,n_1261,n_467,n_185,n_1069,n_465,n_816,n_62,n_1237,n_937,n_276,n_364,n_46,n_888,n_100,n_895,n_1194,n_601,n_803,n_1257,n_978,n_233,n_40,n_271,n_34,n_1227,n_411,n_61,n_537,n_59,n_1157,n_1367,n_451,n_1215,n_641,n_1273,n_1360,n_1083,n_1059,n_1200,n_1259,n_715,n_628,n_181,n_45,n_358,n_788,n_1161,n_908,n_376,n_550,n_899,n_371,n_998,n_814,n_43,n_663,n_42,n_183,n_1153,wire1671,wire1675,wire1306,wire1310,wire1313,wire1318,wire1322,wire1326,wire1330,wire1334,wire1338,wire1342,wire1346,wire1350,wire1354,wire1358,wire1359,wire1360,wire1361,wire1362,wire1363,wire1364,wire1368,wire1372,wire1376,wire1380,wire1384,wire1388,wire1392,wire1396,wire1400,wire1401,wire1402,wire1403,wire1404,wire1405,wire1406,wire1407,wire1408,wire1412,wire1416,wire1420,wire1424,wire1428,wire1432,n_711,n_1290,n_1075,n_725,n_447,n_990,n_168,n_883,n_731,n_1026,n_709,n_994,n_449,n_1322,n_1253,n_1358,n_740,n_1341,n_1114,n_713,n_368,n_515,n_1077,n_1047,n_1151,n_1042,n_267,n_1404,n_1107,n_354,n_1351,n_1268,n_360,n_700,n_548,n_835,n_461,n_187,n_455,n_818,n_191,n_630,n_362,n_1144,n_544,n_808,n_261,n_1332,n_562,n_541,n_257,n_1336,n_1424,n_554,n_166,n_459,n_350,n_751,n_1090,n_79,n_366,n_633,n_621,n_856,n_720,n_443,wire1503,wire1507,n_263,n_1390,n_531,n_810,n_164,n_897,n_981,n_1155,n_259,n_643,n_273,n_1073,n_985,n_635,n_265,n_1003,n_637,n_457,n_348,n_812,n_1096,n_539,n_624,n_1385,n_1081,n_374,n_1128,n_799,n_723,n_1013,n_1310,n_826,n_533,n_734,n_1255,n_282,n_1406,n_1369,n_189,n_893,n_886,n_441,n_278,n_535,n_284,n_1348,n_172,n_453,n_321,n_352,n_1021,n_1338,n_646,n_177,n_1283,n_845,n_626,n_546,n_356,n_170,n_901,n_179,n_1139,n_801,n_1432,n_1300,n_1439,n_445,n_656,n_996,n_1524,n_1525,wire1758,wire1121,wire1301,n_80,wire1314,n_78,n_76,n_75,n_74,n_72,n_71,n_70,n_69,n_68,n_66,n_65,n_98,n_82,n_86,n_83,n_91,n_92,n_57,n_56,n_55,n_54,n_53,n_52,n_51,n_50,n_49,n_97,n_85,n_95,n_84,n_81,n_94,n_96,n_93,n_39,n_38,n_37,n_36,n_33,n_32,n_7,n_6,wire1122,wire1267,wire1269,wire1271,wire1273,wire1275,wire1277,wire1278,wire1280,wire1281,wire1283,wire1284,wire1287,wire1289,wire1291,wire1293,wire1295,wire1296,wire1297,wire1298,wire1299,wire1300,n_122,n_129,n_114,n_131,wire1302,n_135,wire1303,n_141,wire1307,wire1311,n_113,n_133,n_139,wire1312,n_145,n_137,n_99,wire1123,wire1274,wire1276,n_117,wire1279,n_121,wire1282,n_110,n_119,wire1285,wire1288,wire1290,wire1292,wire1294,n_109,n_108,n_106,n_105,n_103,n_102,n_112,n_116,n_120,n_90,n_88,n_118,wire1235,wire1237,wire1245,wire1247,wire1249,wire1258,wire1259,wire1260,wire1262,wire1263,wire1264,wire1266,n_138,n_136,n_132,n_140,wire1286,n_130,n_123,n_115,n_134,n_107,n_104,n_101,wire1233,wire1234,wire1236,wire1238,wire1239,wire1240,wire1241,wire1244,n_143,wire1251,wire1252,wire1253,wire1254,wire1255,wire1256,n_126,n_125,n_124,wire1261,n_155,n_147,n_157,wire1265,n_144,wire1268,wire1270,wire1272,n_128,wire1035,wire1224,n_184,n_186,wire1242,n_182,wire1248,n_149,n_156,n_148,n_154,n_150,n_158,wire1257,n_159,n_151,n_146,n_142,wire1036,wire1185,wire1192,wire1206,wire1219,wire1220,wire1221,n_174,wire1230,wire1232,n_167,n_171,n_180,n_169,n_178,n_165,n_173,n_188,wire1246,n_162,wire1250,n_152,wire1176,wire1178,wire1187,wire1189,wire1190,wire1191,wire1195,wire1208,wire1210,wire1211,wire1216,wire1218,n_196,n_202,n_203,wire1222,wire1223,wire1225,wire1226,wire1227,wire1228,wire1229,wire1231,n_153,wire1243,n_160,n_163,n_208,wire1179,wire1186,wire1193,wire1196,wire1197,wire1205,wire1207,wire1214,n_195,n_194,n_198,n_201,n_199,n_200,n_193,n_197,n_190,n_175,n_192,n_209,wire1149,wire1177,wire1183,wire1188,n_216,n_222,n_226,n_232,wire1194,n_220,n_223,n_236,wire1198,wire1199,wire1200,wire1201,wire1202,wire1203,wire1204,n_227,n_238,wire1209,n_214,n_218,wire1212,wire1213,wire1215,wire1217,wire1756,n_249,n_224,n_215,n_221,n_229,n_219,n_212,n_217,n_225,n_213,n_228,n_206,n_205,n_207,n_211,wire1757,wire1124,wire1150,wire1151,wire1152,wire1153,wire1154,wire1155,wire1156,wire1157,wire1158,wire1166,wire1167,wire1168,wire1169,wire1170,wire1171,wire1172,wire1173,wire1174,n_230,wire1180,wire1181,wire1182,wire1184,n_1566,n_286,wire1142,wire1159,wire1165,n_245,n_241,n_244,n_240,n_243,n_247,n_242,n_248,n_246,wire1175,n_234,n_237,n_231,n_235,wire1077,wire1141,wire1145,wire1146,wire1148,n_274,n_264,n_262,n_272,n_270,n_260,n_266,n_268,n_258,wire1161,wire1162,wire1163,wire1164,n_253,n_239,n_318,wire1107,wire1109,wire1111,wire1112,wire1113,wire1114,wire1116,wire1117,wire1118,wire1131,wire1132,wire1133,wire1134,wire1135,wire1136,wire1137,wire1138,wire1139,n_283,wire1160,n_250,n_252,n_251,n_254,wire1054,wire1093,wire1126,n_291,n_295,n_294,n_290,n_288,n_289,n_292,n_287,n_293,n_279,wire1143,n_277,wire1147,n_285,n_256,n_373,wire1090,wire1091,wire1095,wire1098,wire1099,wire1100,wire1101,wire1102,wire1103,wire1104,wire1105,wire1106,wire1108,wire1110,n_309,n_312,n_303,wire1115,n_311,n_307,n_305,wire1119,wire1125,n_298,wire1127,wire1128,wire1140,wire1144,n_319,wire1037,wire1086,wire1094,n_327,n_313,n_302,n_317,n_310,n_306,n_304,n_308,n_314,n_330,n_324,n_315,n_301,n_297,n_299,n_280,n_275,n_1412,wire1062,wire1063,wire1064,wire1066,wire1067,wire1068,wire1069,wire1079,wire1080,wire1081,wire1082,wire1083,wire1084,wire1085,n_325,wire1087,wire1088,wire1089,n_326,wire1092,n_328,wire1096,wire1097,wire1120,wire1130,wire1754,wire1055,wire1058,wire1072,wire1073,n_333,n_338,n_339,n_335,n_336,n_334,n_340,n_329,n_332,n_323,n_331,n_316,n_296,wire1755,wire1052,wire1057,wire1059,n_349,n_353,n_363,wire1065,n_351,n_361,n_357,n_359,wire1070,wire1071,n_346,n_343,wire1074,wire1078,n_322,n_1565,wire1023,wire1025,wire1026,wire1027,wire1028,wire1030,wire1032,wire1044,wire1045,wire1046,wire1047,wire1049,wire1050,wire1051,n_372,wire1056,n_369,wire1060,n_344,n_347,n_342,wire1075,wire1076,n_337,wire1004,wire1006,wire1038,wire1041,n_378,n_383,n_379,n_380,n_382,n_385,n_381,n_375,n_377,n_367,n_355,n_345,n_341,wire997,wire1008,wire1009,wire1016,wire1017,wire1018,wire1019,wire1020,wire1021,wire1022,n_396,wire1024,n_406,n_398,n_400,wire1029,wire1031,n_408,wire1033,wire1034,n_392,n_391,wire1042,wire1048,wire1053,n_423,wire1061,wire1000,wire1003,wire1005,wire1007,n_407,n_399,n_402,n_403,n_397,n_395,n_405,n_404,n_422,n_393,n_390,n_389,n_384,n_370,n_365,wire975,wire976,wire977,wire979,wire980,wire981,wire990,wire991,wire992,wire994,wire995,wire996,wire998,wire999,n_419,wire1001,wire1002,n_409,n_416,n_420,n_410,wire1010,wire1011,wire1013,wire1015,n_401,wire1040,wire1043,wire971,wire973,wire978,wire984,wire989,n_432,n_425,n_426,wire993,n_433,n_431,n_427,n_421,n_418,n_415,n_417,n_414,n_388,n_386,wire967,wire970,wire972,n_454,n_446,n_444,n_450,n_452,n_442,wire983,n_435,wire985,wire986,n_437,n_430,wire1012,wire1014,wire1752,wire940,wire942,wire943,wire944,wire946,wire948,wire958,wire959,wire960,wire962,wire963,wire964,n_460,n_464,n_448,n_436,n_438,n_439,n_412,n_413,wire1753,wire927,wire931,wire945,wire953,wire955,n_473,n_476,n_470,wire961,n_474,n_475,n_471,n_458,wire968,n_466,n_462,wire974,wire987,wire988,n_1564,wire923,wire925,wire930,wire933,wire934,wire935,wire936,wire937,wire938,wire941,n_487,n_492,n_496,wire947,n_498,wire952,n_477,wire954,n_480,wire956,n_472,wire965,wire982,n_434,n_428,wire918,wire921,wire928,wire932,n_486,n_491,n_495,n_489,n_493,n_497,wire939,n_508,n_488,n_494,n_484,n_478,n_481,wire969,n_456,n_440,wire1750,wire894,wire895,wire896,wire897,wire899,wire900,wire908,wire909,wire910,wire911,wire913,wire914,wire917,n_506,wire919,n_501,wire922,wire924,wire926,n_505,wire929,n_502,n_504,n_500,wire957,wire966,n_521,wire1751,wire887,wire889,wire904,wire906,n_513,n_520,n_514,n_519,n_518,n_517,n_503,n_507,n_510,n_509,n_479,n_468,n_1563,wire888,wire891,wire892,n_534,n_540,n_542,n_532,n_538,n_536,wire902,wire903,n_526,wire905,n_528,wire912,wire915,wire920,n_499,wire950,wire951,wire853,wire861,wire862,wire863,wire865,wire868,wire878,wire879,wire880,wire881,wire883,wire884,n_545,n_553,wire890,n_527,n_523,n_524,wire907,n_512,n_490,n_482,wire844,wire846,wire871,wire875,n_560,n_561,n_556,n_564,n_559,n_558,n_551,n_547,n_555,n_525,n_516,wire916,wire1748,wire842,wire848,wire852,n_585,wire854,wire855,wire856,wire857,wire858,wire859,n_577,n_587,wire864,n_583,wire869,wire870,n_571,wire872,wire874,n_570,wire885,n_549,wire898,n_511,wire1749,wire837,wire841,wire845,wire847,wire851,n_576,n_586,n_582,n_597,n_584,n_580,n_581,n_591,n_565,n_572,wire873,n_569,wire886,n_530,wire901,n_1562,wire812,wire813,wire814,wire815,wire818,wire827,wire828,wire829,wire830,wire832,wire836,n_588,wire838,wire839,n_598,wire843,n_593,n_589,wire849,n_599,n_566,wire876,wire882,n_619,wire893,n_529,wire805,wire807,wire819,wire824,n_606,n_600,n_605,n_608,n_607,n_592,n_594,n_590,wire840,n_595,n_596,n_557,n_563,n_543,wire806,wire808,wire809,wire811,n_629,n_627,n_631,n_625,n_622,n_618,wire820,wire821,wire822,wire823,n_616,wire833,wire834,n_604,wire860,wire867,wire877,wire779,wire781,wire782,wire783,wire785,wire796,wire797,wire798,wire799,wire803,n_634,n_640,n_609,n_617,n_612,n_615,n_575,n_574,n_568,wire755,wire771,wire791,wire794,n_650,n_652,n_651,n_649,n_648,n_642,n_644,n_638,n_636,wire825,wire831,n_603,wire835,wire850,wire763,wire765,wire767,wire773,wire774,wire775,wire776,wire777,wire778,wire780,n_673,n_671,wire784,n_666,wire789,wire790,n_662,wire792,wire793,n_654,wire800,wire816,n_611,n_602,n_578,wire756,wire757,wire762,wire772,n_668,n_672,n_670,n_685,n_665,n_683,n_669,n_653,n_660,n_659,n_658,wire801,n_623,wire817,wire826,wire1746,wire732,wire733,wire734,wire735,wire748,wire749,wire750,wire753,n_681,n_686,wire758,wire759,wire760,wire761,n_676,wire764,wire766,n_684,n_687,n_677,n_647,n_613,n_610,wire1747,wire726,wire727,wire730,wire740,wire741,wire745,n_695,n_694,n_693,wire751,n_692,n_682,n_690,n_680,n_688,n_689,wire786,wire795,wire802,wire810,wire1744,n_1561,wire724,wire725,wire729,n_714,n_710,n_716,n_712,wire739,n_703,n_702,wire742,wire743,n_698,n_667,wire787,n_717,wire804,n_632,wire1745,wire700,wire702,wire704,wire705,wire718,wire719,wire720,wire721,n_728,n_724,n_726,n_699,n_704,n_705,n_691,wire752,n_657,n_645,n_1560,wire684,wire688,wire689,wire710,wire711,wire712,n_739,n_736,n_738,n_737,wire722,n_721,n_732,n_730,wire736,wire746,wire747,n_697,wire768,wire770,wire788,wire675,wire682,wire686,wire696,wire697,wire698,wire699,wire701,wire703,n_759,n_755,wire708,wire709,n_747,n_744,n_745,wire715,n_708,n_674,n_675,n_664,wire676,wire678,wire679,wire685,n_768,wire690,n_758,n_754,n_757,n_769,n_775,n_756,n_750,n_748,n_746,n_735,wire737,wire744,n_701,n_696,wire754,wire647,wire652,wire653,wire654,wire661,wire669,wire670,wire671,wire673,n_767,n_771,wire677,n_778,n_766,wire680,wire681,wire683,n_764,wire687,n_770,wire706,wire713,wire716,wire728,wire731,n_707,n_678,wire644,wire648,wire660,n_787,wire662,n_782,n_781,n_783,n_774,n_773,n_763,n_772,n_753,n_722,n_719,wire738,wire1742,wire642,wire643,wire645,n_811,n_802,n_800,n_804,wire658,wire659,n_786,n_791,wire665,wire672,n_777,n_823,wire714,n_741,n_706,wire1743,wire602,wire616,wire617,wire619,wire633,wire637,wire638,wire639,wire641,n_813,n_817,wire656,n_793,n_792,wire663,n_790,n_785,wire695,wire707,n_743,wire723,n_1559,wire600,wire606,wire628,wire630,n_831,n_820,n_825,n_821,n_819,n_815,n_809,n_794,wire666,wire692,wire693,n_765,wire717,n_733,wire598,n_859,wire608,wire612,wire614,n_840,wire618,wire620,wire622,wire625,wire626,wire627,n_828,wire629,n_833,wire634,n_827,n_784,wire664,n_762,n_752,n_742,wire597,wire601,wire605,wire607,n_864,wire615,n_842,n_849,wire621,n_839,n_858,n_841,n_829,n_832,n_830,wire635,wire649,wire657,n_796,wire667,wire674,wire694,wire569,wire574,wire575,wire581,wire595,wire596,wire599,n_861,n_850,n_853,wire609,wire610,wire611,wire613,n_851,n_860,n_838,n_807,n_789,n_776,n_761,wire563,wire566,wire580,n_871,wire585,wire594,n_866,n_867,n_863,n_855,n_854,n_848,n_852,wire631,n_836,wire646,wire650,wire655,n_795,wire668,wire559,wire564,wire565,wire568,wire570,n_887,n_889,wire578,n_878,wire583,wire584,n_875,wire586,wire588,n_873,wire603,wire624,wire640,n_797,n_806,n_779,wire536,wire538,wire557,wire558,n_904,n_898,n_896,n_885,n_876,n_877,n_872,n_847,wire632,n_822,wire651,wire1738,wire1740,wire521,wire525,wire532,wire546,wire549,wire550,n_911,n_912,wire560,n_894,n_900,n_902,wire587,n_874,n_846,n_916,n_805,wire1739,wire1741,wire514,wire523,wire527,wire534,wire535,wire537,wire539,n_925,wire547,wire548,n_915,n_913,wire551,wire552,n_909,wire567,wire576,n_882,wire589,wire604,wire636,n_1557,n_1558,wire507,wire516,wire517,wire522,wire526,wire533,n_943,n_935,n_934,n_952,wire542,n_921,n_926,n_922,n_892,wire579,n_865,wire591,wire592,wire623,n_834,wire1734,wire487,wire506,wire515,n_939,n_948,wire518,wire519,wire520,n_946,wire524,n_944,n_940,n_947,n_923,wire553,n_881,wire577,n_862,n_857,n_843,wire1735,wire477,wire480,wire485,wire497,wire499,wire502,n_953,wire508,n_951,n_945,n_950,n_949,wire543,n_920,wire562,wire572,n_891,n_884,wire582,wire593,wire1732,n_1555,wire478,wire479,wire481,wire488,wire495,wire496,n_973,wire498,n_964,wire500,n_970,n_961,wire528,wire540,wire561,n_907,n_870,n_869,wire1726,wire1733,wire472,n_999,n_986,n_991,n_982,wire489,n_971,n_969,n_972,n_932,wire544,wire555,n_910,wire571,n_890,wire573,n_1554,wire444,wire447,wire451,wire455,wire461,wire465,wire467,wire471,n_995,n_997,n_993,n_980,wire501,wire529,n_1018,wire541,n_931,wire554,n_906,n_879,wire1730,wire436,wire449,wire452,n_1012,wire462,wire463,wire464,n_1010,n_1015,n_1005,n_1004,wire490,n_965,wire509,n_929,n_918,wire556,wire1731,wire1736,wire432,wire438,wire442,wire443,wire445,wire448,n_1036,n_1040,wire456,n_1009,n_1011,n_1016,wire466,wire482,wire493,n_941,wire511,wire530,n_905,wire1727,n_1553,wire1737,wire437,n_1037,wire439,wire440,wire441,n_1045,n_1031,n_1038,n_1030,wire450,n_1032,n_1023,n_987,wire491,n_955,wire512,n_938,wire545,n_1551,wire1728,n_1556,wire402,wire405,wire406,wire420,wire421,wire423,wire431,n_1046,n_1034,n_1039,n_1029,n_1033,n_1014,wire483,n_975,wire494,wire503,wire504,wire531,n_928,wire1729,wire396,wire401,wire403,wire404,wire414,wire419,n_1054,n_1053,wire422,n_1057,wire424,wire426,n_1051,wire446,wire458,wire474,n_979,n_958,wire513,n_936,n_1552,n_1076,n_1084,n_1078,n_1064,n_1058,n_1056,n_1055,n_1028,wire459,wire473,n_1000,wire484,wire505,n_957,wire1724,wire370,wire372,wire378,wire385,wire388,wire389,n_1091,n_1082,n_1080,n_1074,wire425,n_1052,n_1022,n_988,wire475,n_983,wire492,n_963,wire1725,wire355,wire365,wire366,wire368,wire380,n_1092,wire386,wire387,n_1098,n_1099,wire390,wire395,wire407,wire415,n_1063,wire433,wire453,wire460,wire468,wire469,wire486,n_967,wire1718,n_1550,wire359,wire362,wire364,wire371,n_1125,wire379,n_1109,n_1103,n_1100,n_1102,n_1065,n_1044,n_1110,n_1008,wire476,n_976,wire1719,wire1722,wire354,n_1132,n_1118,wire360,wire361,n_1131,wire363,n_1121,n_1119,wire367,wire369,n_1120,n_1117,n_1097,wire413,n_1062,n_1027,wire470,n_1001,n_1547,wire1720,wire1723,wire317,wire331,wire332,wire337,wire346,wire347,wire350,n_1141,n_1123,n_1124,n_1116,n_1122,wire373,wire381,wire397,wire409,wire410,n_1068,wire427,wire429,wire434,wire457,n_1006,wire1721,n_1549,wire333,wire334,wire335,n_1150,wire344,wire345,n_1136,n_1137,wire348,n_1113,n_1089,n_1050,n_1049,wire430,wire454,n_1020,n_1548,wire318,n_1156,n_1154,n_1133,n_1134,n_1135,n_1142,wire351,n_1108,wire408,n_1067,wire411,wire417,n_1043,wire435,n_1024,wire289,wire296,wire308,wire314,wire315,n_1169,wire327,n_1152,n_1160,wire336,wire339,n_1149,wire356,wire376,wire392,wire399,n_1086,n_1070,wire416,n_1048,n_1041,wire272,wire279,wire291,wire304,wire312,n_1181,n_1183,wire316,n_1164,n_1158,n_1130,wire374,wire391,n_1095,wire394,wire412,n_1061,wire418,wire285,wire288,wire290,wire294,wire297,n_1184,wire309,n_1187,wire313,n_1182,wire338,n_1148,n_1115,n_1087,wire398,n_1085,n_1066,n_1060,wire273,wire280,wire284,n_1206,n_1208,n_1203,wire292,wire293,n_1209,wire301,n_1180,n_1172,wire319,wire325,n_1166,wire349,wire357,wire375,wire382,wire384,wire393,n_1093,n_1094,wire400,wire1708,wire1714,wire244,wire265,wire267,n_1222,n_1213,n_1214,n_1202,wire295,wire298,n_1174,n_1143,wire352,n_1219,wire377,n_1106,n_1105,n_1071,wire1709,wire1710,wire1715,wire240,wire241,wire261,n_1224,wire269,n_1207,n_1196,wire302,n_1165,wire326,n_1129,n_1112,wire383,n_1542,wire1711,n_1545,wire1716,wire245,wire246,n_1235,wire266,wire268,n_1236,wire286,n_1195,wire307,wire321,wire322,n_1178,wire340,wire342,n_1140,n_1104,wire1698,wire1704,n_1543,wire1717,wire235,n_1254,n_1260,n_1256,wire256,wire259,n_1233,n_1230,wire274,n_1186,wire310,wire328,n_1147,n_1146,wire343,wire358,wire1705,n_1546,wire203,wire204,wire209,wire222,wire224,wire225,wire226,wire247,wire250,n_1243,n_1204,wire287,wire320,n_1177,wire323,n_1163,wire329,wire353,n_1126,n_1540,n_1277,n_1282,n_1281,n_1269,n_1258,n_1252,wire260,wire277,n_1201,wire299,wire306,n_1188,n_1189,n_1176,n_1145,n_1138,wire1702,wire194,wire202,n_1303,wire205,wire206,wire208,wire210,wire216,wire223,n_1284,wire248,n_1242,wire263,wire270,wire275,wire281,n_1193,wire300,wire305,n_1199,wire324,wire330,wire1699,wire1703,wire184,wire201,n_1298,n_1299,n_1302,n_1292,wire217,n_1270,wire236,n_1217,wire278,n_1210,n_1191,n_1167,n_1162,n_1537,n_1539,wire173,wire175,wire186,wire190,n_1306,wire195,n_1304,wire207,n_1267,wire249,wire264,wire276,n_1216,wire282,wire303,n_1198,wire311,wire1688,wire1700,wire1706,n_1314,wire185,n_1316,n_1317,n_1313,n_1294,n_1291,wire238,n_1247,wire254,wire258,n_1228,wire271,n_1318,n_1212,n_1170,wire1689,wire1701,wire1707,wire159,wire174,n_1337,wire176,wire177,wire179,n_1324,wire193,wire196,wire215,wire227,wire231,wire251,n_1231,n_1223,wire283,n_1532,n_1538,n_1541,wire1712,wire134,wire156,wire165,n_1328,n_1334,wire183,n_1315,n_1312,wire229,n_1272,wire239,n_1239,wire253,wire255,n_1211,wire1696,wire1713,n_1363,n_1359,n_1339,wire178,n_1325,n_1327,n_1301,wire228,n_1266,wire242,n_1249,n_1238,wire262,wire1682,wire1694,wire1697,n_1544,wire1759,wire116,wire133,wire135,wire137,wire140,wire148,wire155,n_1349,wire167,wire169,n_1344,wire187,wire198,wire218,wire220,n_1275,wire230,wire233,wire237,wire257,n_1234,wire1683,wire1695,n_1536,n_1567,wire126,n_1388,n_1378,n_1380,wire149,n_1357,n_1350,n_1321,wire192,wire213,n_1285,n_1274,n_1250,wire243,n_1244,n_1529,n_1535,n_1399,wire117,wire120,wire127,n_1379,wire141,n_1370,n_1373,n_1343,wire170,wire188,n_1311,n_1295,wire214,wire221,wire234,n_1246,wire1692,wire99,wire104,wire118,n_1408,wire121,wire124,n_1394,n_1387,wire129,wire138,n_1393,wire153,wire161,n_1347,wire180,n_1323,wire211,n_1288,n_1286,wire232,n_1262,wire1693,wire84,wire94,wire106,wire112,n_1413,n_1403,n_1398,n_1392,wire151,n_1362,wire168,n_1331,wire182,wire189,wire197,wire199,wire219,n_1263,wire1684,n_1534,wire83,wire89,wire90,n_1422,wire102,n_1409,n_1410,wire109,n_1421,n_1386,n_1346,wire162,n_1345,n_1417,n_1307,wire212,n_1279,wire1685,wire1690,wire64,wire74,wire80,wire85,wire91,n_1456,wire95,wire98,n_1419,n_1428,wire113,wire128,wire150,n_1355,wire152,n_1356,n_1333,wire200,n_1296,n_1530,wire1686,wire1691,n_1436,n_1470,wire92,n_1429,n_1397,wire122,wire142,wire143,wire145,n_1371,n_1366,wire160,wire164,wire171,wire191,n_1308,wire1687,n_1533,wire67,n_1479,n_1427,wire103,n_1391,n_1377,n_1353,n_1354,wire166,wire181,n_1320,n_1531,wire62,n_1457,wire75,wire88,n_1431,wire110,n_1405,wire144,n_1365,wire146,wire157,n_1342,wire172,n_1326,wire42,wire52,n_1443,wire76,wire97,n_1415,wire111,wire131,wire136,n_1368,n_1382,wire154,n_1352,n_1335,n_1464,n_1483,wire87,n_1430,n_1426,wire107,wire125,wire130,n_1389,wire147,n_1364,wire158,wire44,wire55,wire73,n_1438,wire77,n_1437,n_1407,n_1383,wire132,n_1381,n_1374,n_1361,n_1471,wire50,wire66,wire71,n_1450,n_1447,wire96,wire101,wire108,wire114,wire119,wire123,n_1395,n_1396,wire139,wire1678,wire34,wire39,n_1487,n_1458,wire93,n_1434,wire105,n_1473,n_1400,n_1402,n_1375,wire1679,n_1477,n_1491,wire70,n_1446,n_1425,n_1411,wire115,n_1527,wire1680,wire33,wire46,wire58,wire60,wire63,n_1452,wire78,wire82,n_1433,n_1401,wire1681,n_1480,wire56,n_1461,wire72,n_1444,wire79,n_1442,wire100,n_1528,wire31,wire32,n_1495,n_1451,wire61,n_1519,wire68,n_1445,wire86,n_1423,n_1481,wire43,wire54,n_1459,wire59,n_1460,n_1440,n_1435,wire30,wire40,wire49,wire51,n_1465,n_1463,wire65,wire69,n_1484,n_1499,n_1469,n_1453,n_1449,wire28,wire29,n_1503,wire47,n_1462,wire53,wire57,n_1485,wire38,wire45,n_1468,n_1454,wire27,n_1472,wire48,wire1676,n_1488,n_1507,n_1467,wire1677,wire24,wire26,wire36,wire41,n_1526,n_1489,wire35,wire37,n_1475,wire25,n_1511,n_1476,n_1492,n_1515,wire21,wire23,n_1493,wire22,n_1496,wire18,wire20,n_1497,wire19,n_1500,wire16,wire17,n_1501,wire15,n_1504,wire12,wire14,n_1505,wire13,n_1508,wire10,wire11,n_1509,wire9,n_1512,wire6,wire8,n_1513,wire7,n_1516,wire3,wire5,n_1517,wire4,n_1520,wire1,wire2,n_1521,wire0;

and AND2_1 (wire81, n256, n528);
and AND2_2 (wire163, n256, n511);
and AND2_3 (wire252, n256, n494);
and AND2_4 (wire341, n256, n477);
and AND2_5 (wire428, n256, n460);
and AND2_6 (wire510, n256, n443);
and AND2_7 (wire590, n256, n426);
and AND2_8 (wire691, n256, n409);
and AND2_9 (wire769, n256, n392);
and AND2_10 (wire866, n256, n375);
and AND2_11 (wire949, n256, n358);
and AND2_12 (wire1039, n256, n341);
and AND2_13 (wire1129, n256, n324);
not NOT1_14 (wire1315, keyinput28);
not NOT1_15 (wire1319, keyinput21);
not NOT1_16 (wire1323, keyinput12);
and AND2_17 (wire1325, keyinput12, n154);
not NOT1_18 (wire1327, keyinput29);
not NOT1_19 (wire1331, keyinput6);
not NOT1_20 (wire1335, keyinput14);
not NOT1_21 (wire1339, keyinput18);
not NOT1_22 (wire1343, keyinput5);
not NOT1_23 (wire1347, keyinput1);
not NOT1_24 (wire1351, keyinput15);
and AND2_25 (wire1353, keyinput15, n392);
not NOT1_26 (wire1355, keyinput3);
not NOT1_27 (wire1365, keyinput10);
not NOT1_28 (wire1369, keyinput27);
and AND2_29 (wire1371, keyinput27, n494);
not NOT1_30 (wire1373, keyinput26);
and AND2_31 (wire1375, keyinput26, n35);
not NOT1_32 (wire1377, keyinput23);
not NOT1_33 (wire1381, keyinput31);
not NOT1_34 (wire1385, keyinput22);
not NOT1_35 (wire1389, keyinput19);
not NOT1_36 (wire1393, keyinput11);
not NOT1_37 (wire1397, keyinput25);
or OR2_38 (wire1409, n86, keyinput20);
and AND2_39 (wire1410, n86, keyinput20);
or OR2_40 (wire1413, n188, keyinput8);
and AND2_41 (wire1414, n188, keyinput8);
or OR2_42 (wire1417, n528, keyinput30);
and AND2_43 (wire1418, n528, keyinput30);
or OR2_44 (wire1421, n341, keyinput9);
and AND2_45 (wire1422, n341, keyinput9);
or OR2_46 (wire1425, n120, keyinput16);
and AND2_47 (wire1426, n120, keyinput16);
or OR2_48 (wire1429, n409, keyinput17);
and AND2_49 (wire1430, n409, keyinput17);
or OR2_50 (wire1500, n324, keyinput7);
and AND2_51 (wire1501, n324, keyinput7);
or OR2_52 (wire1504, n239, keyinput2);
and AND2_53 (wire1505, n239, keyinput2);
and AND2_54 (wire1578, n188, n290);
and AND2_55 (wire1579, n35, n392);
and AND2_56 (wire1580, n120, n290);
and AND2_57 (wire1581, n86, n494);
and AND2_58 (wire1582, n1, n494);
and AND2_59 (wire1583, n1, n409);
and AND2_60 (wire1584, n86, n290);
and AND2_61 (wire1585, n239, n307);
and AND2_62 (wire1586, n35, n443);
and AND2_63 (wire1587, n222, n324);
and AND2_64 (wire1588, n137, n290);
and AND2_65 (wire1589, n35, n409);
and AND2_66 (wire1590, n222, n426);
and AND2_67 (wire1591, n35, n375);
and AND2_68 (wire1592, n35, n358);
and AND2_69 (wire1593, n1, n477);
and AND2_70 (wire1594, n35, n324);
and AND2_71 (wire1595, n222, n375);
and AND2_72 (wire1596, n222, n409);
and AND2_73 (wire1597, n35, n290);
and AND2_74 (wire1598, n205, n443);
and AND2_75 (wire1599, n239, n494);
and AND2_76 (wire1600, n222, n443);
and AND2_77 (wire1601, n103, n494);
and AND2_78 (wire1602, n222, n307);
and AND2_79 (wire1603, n1, n460);
and AND2_80 (wire1604, n205, n290);
and AND2_81 (wire1605, n154, n443);
and AND2_82 (wire1606, n171, n443);
and AND2_83 (wire1607, n205, n494);
and AND2_84 (wire1608, n222, n528);
and AND2_85 (wire1609, n222, n494);
and AND2_86 (wire1610, n222, n358);
and AND2_87 (wire1611, n86, n307);
and AND2_88 (wire1612, n239, n477);
and AND2_89 (wire1613, n1, n358);
and AND2_90 (wire1614, n35, n426);
and AND2_91 (wire1615, n69, n290);
and AND2_92 (wire1616, n188, n494);
and AND2_93 (wire1617, n188, n443);
and AND2_94 (wire1618, n1, n324);
and AND2_95 (wire1619, n222, n341);
and AND2_96 (wire1620, n52, n290);
and AND2_97 (wire1621, n86, n443);
and AND2_98 (wire1622, n256, n273);
and AND2_99 (wire1623, n120, n443);
and AND2_100 (wire1624, n120, n494);
and AND2_101 (wire1625, n239, n392);
and AND2_102 (wire1626, n86, n426);
and AND2_103 (wire1627, n52, n511);
and AND2_104 (wire1628, n239, n460);
and AND2_105 (wire1629, n239, n324);
and AND2_106 (wire1630, n103, n290);
and AND2_107 (wire1631, n86, n324);
and AND2_108 (wire1632, n1, n528);
and AND2_109 (wire1633, n171, n494);
and AND2_110 (wire1634, n239, n358);
and AND2_111 (wire1635, n222, n290);
and AND2_112 (wire1636, n86, n375);
and AND2_113 (wire1637, n18, n290);
and AND2_114 (wire1638, n69, n494);
and AND2_115 (wire1639, n239, n528);
and AND2_116 (wire1640, n86, n358);
and AND2_117 (wire1641, n154, n494);
and AND2_118 (wire1642, n1, n392);
and AND2_119 (wire1643, n239, n511);
and AND2_120 (wire1644, n222, n511);
and AND2_121 (wire1645, n35, n477);
and AND2_122 (wire1646, n222, n460);
and AND2_123 (wire1647, n137, n494);
and AND2_124 (wire1648, n1, n511);
and AND2_125 (wire1649, n86, n409);
and AND2_126 (wire1650, n86, n392);
and AND2_127 (wire1651, n35, n307);
and AND2_128 (wire1652, n154, n290);
and AND2_129 (wire1653, n86, n341);
and AND2_130 (wire1654, n239, n426);
and AND2_131 (wire1655, n222, n477);
and AND2_132 (wire1656, n137, n443);
and AND2_133 (wire1657, n1, n341);
and AND2_134 (wire1658, n1, n375);
and AND2_135 (wire1659, n1, n443);
and AND2_136 (wire1660, n35, n341);
and AND2_137 (wire1661, n35, n460);
and AND2_138 (wire1662, n1, n426);
and AND2_139 (wire1663, n171, n290);
and AND2_140 (wire1664, n222, n392);
and AND2_141 (wire1665, n1, n290);
and AND2_142 (wire1666, n1, n307);
and AND2_143 (wire1667, n35, n494);
not NOT1_144 (n_67, n290);
not NOT1_145 (n_4, n35);
not NOT1_146 (n_5, n86);
not NOT1_147 (n_29, n409);
not NOT1_148 (n_12, n426);
not NOT1_149 (n_13, n341);
not NOT1_150 (n_15, n324);
not NOT1_151 (n_26, n460);
not NOT1_152 (n_21, n171);
not NOT1_153 (n_27, n188);
not NOT1_154 (n_73, n511);
not NOT1_155 (n_19, n154);
not NOT1_156 (n_20, n137);
not NOT1_157 (n_22, n69);
not NOT1_158 (n_31, n103);
not NOT1_159 (n_1, keyinput24);
not NOT1_160 (n_0, keyinput13);
not NOT1_161 (n_8, n273);
not NOT1_162 (n_9, n1);
not NOT1_163 (n_16, n494);
not NOT1_164 (n_23, n239);
not NOT1_165 (n_24, n443);
not NOT1_166 (n_25, n307);
not NOT1_167 (n_28, n358);
not NOT1_168 (n_11, n392);
not NOT1_169 (n_14, n528);
not NOT1_170 (n_30, n477);
not NOT1_171 (n_17, n205);
not NOT1_172 (n_89, n375);
not NOT1_173 (n_18, n120);
not NOT1_174 (n_87, n52);
not NOT1_175 (n_77, n18);
not NOT1_176 (wire1668, n256);
not NOT1_177 (wire1669, keyinput0);
and AND2_178 (wire1670, n256, keyinput0);
not NOT1_179 (wire1672, n222);
not NOT1_180 (wire1673, keyinput4);
and AND2_181 (wire1674, n222, keyinput4);
or OR2_182 (wire1304, n375, n_0);
or OR2_183 (wire1305, n_89, keyinput13);
or OR2_184 (wire1308, n52, n_1);
or OR2_185 (wire1309, n_87, keyinput24);
and AND2_186 (wire1316, wire1315, n18);
and AND2_187 (wire1317, keyinput28, n_77);
and AND2_188 (wire1320, wire1319, n443);
and AND2_189 (wire1321, keyinput21, n_24);
and AND2_190 (wire1324, wire1323, n_19);
and AND2_191 (wire1328, wire1327, n511);
and AND2_192 (wire1329, keyinput29, n_73);
and AND2_193 (wire1332, wire1331, n205);
and AND2_194 (wire1333, keyinput6, n_17);
and AND2_195 (wire1336, wire1335, n137);
and AND2_196 (wire1337, keyinput14, n_20);
and AND2_197 (wire1340, wire1339, n103);
and AND2_198 (wire1341, keyinput18, n_31);
and AND2_199 (wire1344, wire1343, n273);
and AND2_200 (wire1345, keyinput5, n_8);
and AND2_201 (wire1348, wire1347, n290);
and AND2_202 (wire1349, keyinput1, n_67);
and AND2_203 (wire1352, wire1351, n_11);
and AND2_204 (wire1356, wire1355, n307);
and AND2_205 (wire1357, keyinput3, n_25);
and AND2_206 (wire1366, wire1365, n171);
and AND2_207 (wire1367, keyinput10, n_21);
and AND2_208 (wire1370, wire1369, n_16);
and AND2_209 (wire1374, wire1373, n_4);
and AND2_210 (wire1378, wire1377, n460);
and AND2_211 (wire1379, keyinput23, n_26);
and AND2_212 (wire1382, wire1381, n1);
and AND2_213 (wire1383, keyinput31, n_9);
and AND2_214 (wire1386, wire1385, n69);
and AND2_215 (wire1387, keyinput22, n_22);
and AND2_216 (wire1390, wire1389, n426);
and AND2_217 (wire1391, keyinput19, n_12);
and AND2_218 (wire1394, wire1393, n358);
and AND2_219 (wire1395, keyinput11, n_28);
and AND2_220 (wire1398, wire1397, n477);
and AND2_221 (wire1399, keyinput25, n_30);
not NOT1_222 (wire1411, wire1410);
not NOT1_223 (wire1415, wire1414);
not NOT1_224 (wire1419, wire1418);
not NOT1_225 (wire1423, wire1422);
not NOT1_226 (wire1427, wire1426);
not NOT1_227 (wire1431, wire1430);
or OR2_228 (wire1433, n_31, n_29);
or OR2_229 (wire1434, n_31, n_73);
or OR2_230 (wire1435, n_87, n_30);
or OR2_231 (wire1436, n_87, n_29);
or OR2_232 (wire1437, n_28, n_27);
or OR2_233 (wire1438, n_31, n_26);
or OR2_234 (wire1439, n_25, n_87);
or OR2_235 (wire1440, n_24, n_23);
or OR2_236 (wire1441, n_22, n_29);
or OR2_237 (wire1442, n_21, n_26);
or OR2_238 (wire1443, n_20, n_29);
or OR2_239 (wire1444, n_77, n_26);
or OR2_240 (wire1445, n_28, n_19);
or OR2_241 (wire1446, n_19, n_73);
or OR2_242 (wire1447, n_77, n_73);
or OR2_243 (wire1448, n_22, n_14);
or OR2_244 (wire1449, n_29, n_27);
or OR2_245 (wire1450, n_27, n_73);
or OR2_246 (wire1451, n_19, n_30);
or OR2_247 (wire1452, n_18, n_29);
or OR2_248 (wire1453, n_13, n_87);
or OR2_249 (wire1454, n_89, n_23);
or OR2_250 (wire1455, n_5, n_30);
or OR2_251 (wire1456, n_17, n_26);
or OR2_252 (wire1457, n_77, n_16);
or OR2_253 (wire1458, n_27, n_26);
or OR2_254 (wire1459, n_15, n_31);
or OR2_255 (wire1460, n_20, n_14);
or OR2_256 (wire1461, n_20, n_30);
or OR2_257 (wire1462, n_13, n_17);
or OR2_258 (wire1463, n_17, n_73);
or OR2_259 (wire1464, n_22, n_73);
or OR2_260 (wire1465, n_13, n_18);
or OR2_261 (wire1466, n_29, n_23);
or OR2_262 (wire1467, n_89, n_27);
or OR2_263 (wire1468, n_12, n_21);
or OR2_264 (wire1469, n_28, n_22);
or OR2_265 (wire1470, n_25, n_31);
or OR2_266 (wire1471, n_28, n_17);
or OR2_267 (wire1472, n_22, n_12);
or OR2_268 (wire1473, n_25, n_22);
or OR2_269 (wire1474, n_19, n_11);
or OR2_270 (wire1475, n_13, n_27);
or OR2_271 (wire1476, n_30, n_17);
or OR2_272 (wire1477, n_89, n_87);
or OR2_273 (wire1478, n_77, n_12);
or OR2_274 (wire1479, n_15, n_17);
or OR2_275 (wire1480, n_21, n_73);
or OR2_276 (wire1481, n_89, n_17);
or OR2_277 (wire1482, n_89, n_21);
or OR2_278 (wire1483, n_15, n_20);
or OR2_279 (wire1484, n_77, n_14);
or OR2_280 (wire1485, n_21, n_14);
or OR2_281 (wire1486, n_89, n_22);
or OR2_282 (wire1487, n_25, n_27);
or OR2_283 (wire1488, n_28, n_87);
or OR2_284 (wire1489, n_13, n_21);
or OR2_285 (wire1490, n_29, n_17);
or OR2_286 (wire1491, n_31, n_30);
or OR2_287 (wire1492, n_67, n_23);
or OR2_288 (wire1493, n_13, n_77);
or OR2_289 (wire1494, n_87, n_11);
or OR2_290 (wire1495, n_18, n_11);
or OR2_291 (wire1496, n_12, n_17);
or OR2_292 (wire1497, n_77, n_29);
or OR2_293 (wire1498, n_28, n_20);
or OR2_294 (wire1499, n_9, n_8);
not NOT1_295 (wire1502, wire1501);
not NOT1_296 (wire1506, wire1505);
or OR2_297 (wire1508, n_15, n_21);
or OR2_298 (wire1509, n_18, n_14);
or OR2_299 (wire1510, n_89, n_18);
or OR2_300 (wire1511, n_20, n_12);
or OR2_301 (wire1512, n_25, n_19);
or OR2_302 (wire1513, n_87, n_24);
or OR2_303 (wire1514, n_5, n_26);
or OR2_304 (wire1515, n_87, n_16);
or OR2_305 (wire1516, n_15, n_18);
or OR2_306 (wire1517, n_22, n_11);
or OR2_307 (wire1518, n_15, n_19);
or OR2_308 (wire1519, n_77, n_30);
or OR2_309 (wire1520, n_87, n_26);
or OR2_310 (wire1521, n_21, n_11);
or OR2_311 (wire1522, n_15, n_27);
or OR2_312 (wire1523, n_18, n_26);
or OR2_313 (wire1524, n_77, n_11);
or OR2_314 (wire1525, n_28, n_77);
or OR2_315 (wire1526, n_13, n_20);
or OR2_316 (wire1527, n_87, n_12);
or OR2_317 (wire1528, n_18, n_30);
or OR2_318 (wire1529, n_89, n_19);
or OR2_319 (wire1530, n_31, n_11);
or OR2_320 (wire1531, n_31, n_14);
or OR2_321 (wire1532, n_22, n_30);
or OR2_322 (wire1533, n_13, n_22);
or OR2_323 (wire1534, n_21, n_30);
or OR2_324 (wire1535, n_18, n_12);
or OR2_325 (wire1536, n_19, n_29);
or OR2_326 (wire1537, n_20, n_26);
or OR2_327 (wire1538, n_20, n_73);
or OR2_328 (wire1539, n_19, n_12);
or OR2_329 (wire1540, n_89, n_31);
or OR2_330 (wire1541, n_29, n_21);
or OR2_331 (wire1542, n_4, n_73);
or OR2_332 (wire1543, n_15, n_87);
or OR2_333 (wire1544, n_19, n_14);
or OR2_334 (wire1545, n_5, n_14);
or OR2_335 (wire1546, n_25, n_77);
or OR2_336 (wire1547, n_77, n_24);
or OR2_337 (wire1548, n_31, n_24);
or OR2_338 (wire1549, n_28, n_31);
or OR2_339 (wire1550, n_15, n_77);
or OR2_340 (wire1551, n_89, n_20);
or OR2_341 (wire1552, n_15, n_22);
or OR2_342 (wire1553, n_87, n_14);
or OR2_343 (wire1554, n_25, n_20);
or OR2_344 (wire1555, n_28, n_18);
or OR2_345 (wire1556, n_13, n_23);
or OR2_346 (wire1557, n_13, n_19);
or OR2_347 (wire1558, n_19, n_26);
or OR2_348 (wire1559, n_4, n_14);
or OR2_349 (wire1560, n_11, n_27);
or OR2_350 (wire1561, n_25, n_17);
or OR2_351 (wire1562, n_5, n_73);
or OR2_352 (wire1563, n_12, n_27);
or OR2_353 (wire1564, n_20, n_11);
or OR2_354 (wire1565, n_89, n_77);
or OR2_355 (wire1566, n_13, n_31);
or OR2_356 (wire1567, n_25, n_18);
or OR2_357 (wire1568, n_22, n_24);
or OR2_358 (wire1569, n_25, n_21);
or OR2_359 (wire1570, n_27, n_30);
or OR2_360 (wire1571, n_31, n_12);
or OR2_361 (wire1572, n_27, n_14);
or OR2_362 (wire1573, n_18, n_73);
or OR2_363 (wire1574, n_17, n_14);
or OR2_364 (wire1575, n_28, n_21);
or OR2_365 (wire1576, n_11, n_17);
or OR2_366 (wire1577, n_22, n_26);
not NOT1_367 (n_63, wire1578);
not NOT1_368 (n_639, wire1579);
not NOT1_369 (n_47, wire1580);
not NOT1_370 (n_1168, wire1581);
not NOT1_371 (n_1159, wire1582);
not NOT1_372 (n_729, wire1583);
not NOT1_373 (n_58, wire1584);
not NOT1_374 (n_127, wire1585);
not NOT1_375 (n_903, wire1586);
not NOT1_376 (n_255, wire1587);
not NOT1_377 (n_44, wire1588);
not NOT1_378 (n_727, wire1589);
not NOT1_379 (n_868, wire1590);
not NOT1_380 (n_552, wire1591);
not NOT1_381 (n_463, wire1592);
not NOT1_382 (n_1079, wire1593);
not NOT1_383 (n_269, wire1594);
not NOT1_384 (n_567, wire1595);
not NOT1_385 (n_760, wire1596);
not NOT1_386 (n_60, wire1597);
not NOT1_387 (n_956, wire1598);
not NOT1_388 (n_1175, wire1599);
not NOT1_389 (n_962, wire1600);
not NOT1_390 (n_1179, wire1601);
not NOT1_391 (n_161, wire1602);
not NOT1_392 (n_992, wire1603);
not NOT1_393 (n_41, wire1604);
not NOT1_394 (n_919, wire1605);
not NOT1_395 (n_930, wire1606);
not NOT1_396 (n_1245, wire1607);
not NOT1_397 (n_1448, wire1608);
not NOT1_398 (n_1261, wire1609);
not NOT1_399 (n_467, wire1610);
not NOT1_400 (n_185, wire1611);
not NOT1_401 (n_1069, wire1612);
not NOT1_402 (n_465, wire1613);
not NOT1_403 (n_816, wire1614);
not NOT1_404 (n_62, wire1615);
not NOT1_405 (n_1237, wire1616);
not NOT1_406 (n_937, wire1617);
not NOT1_407 (n_276, wire1618);
not NOT1_408 (n_364, wire1619);
not NOT1_409 (n_46, wire1620);
not NOT1_410 (n_888, wire1621);
not NOT1_411 (n_100, wire1622);
not NOT1_412 (n_895, wire1623);
not NOT1_413 (n_1194, wire1624);
not NOT1_414 (n_601, wire1625);
not NOT1_415 (n_803, wire1626);
not NOT1_416 (n_1257, wire1627);
not NOT1_417 (n_978, wire1628);
not NOT1_418 (n_233, wire1629);
not NOT1_419 (n_40, wire1630);
not NOT1_420 (n_271, wire1631);
not NOT1_421 (n_34, wire1632);
not NOT1_422 (n_1227, wire1633);
not NOT1_423 (n_411, wire1634);
not NOT1_424 (n_61, wire1635);
not NOT1_425 (n_537, wire1636);
not NOT1_426 (n_59, wire1637);
not NOT1_427 (n_1157, wire1638);
not NOT1_428 (n_1367, wire1639);
not NOT1_429 (n_451, wire1640);
not NOT1_430 (n_1215, wire1641);
not NOT1_431 (n_641, wire1642);
not NOT1_432 (n_1273, wire1643);
not NOT1_433 (n_1360, wire1644);
not NOT1_434 (n_1083, wire1645);
not NOT1_435 (n_1059, wire1646);
not NOT1_436 (n_1200, wire1647);
not NOT1_437 (n_1259, wire1648);
not NOT1_438 (n_715, wire1649);
not NOT1_439 (n_628, wire1650);
not NOT1_440 (n_181, wire1651);
not NOT1_441 (n_45, wire1652);
not NOT1_442 (n_358, wire1653);
not NOT1_443 (n_788, wire1654);
not NOT1_444 (n_1161, wire1655);
not NOT1_445 (n_908, wire1656);
not NOT1_446 (n_376, wire1657);
not NOT1_447 (n_550, wire1658);
not NOT1_448 (n_899, wire1659);
not NOT1_449 (n_371, wire1660);
not NOT1_450 (n_998, wire1661);
not NOT1_451 (n_814, wire1662);
not NOT1_452 (n_43, wire1663);
not NOT1_453 (n_663, wire1664);
not NOT1_454 (n_42, wire1665);
not NOT1_455 (n_183, wire1666);
not NOT1_456 (n_1153, wire1667);
and AND2_457 (wire1671, wire1668, wire1669);
and AND2_458 (wire1675, wire1672, wire1673);
and AND2_459 (wire1306, wire1305, wire1304);
and AND2_460 (wire1310, wire1309, wire1308);
or OR4_461 (wire1313, n_100, n528, n171, n1);
or OR2_462 (wire1318, wire1317, wire1316);
or OR2_463 (wire1322, wire1321, wire1320);
or OR2_464 (wire1326, wire1325, wire1324);
or OR2_465 (wire1330, wire1329, wire1328);
or OR2_466 (wire1334, wire1333, wire1332);
or OR2_467 (wire1338, wire1337, wire1336);
or OR2_468 (wire1342, wire1341, wire1340);
or OR2_469 (wire1346, wire1345, wire1344);
or OR2_470 (wire1350, wire1349, wire1348);
or OR2_471 (wire1354, wire1353, wire1352);
or OR2_472 (wire1358, wire1357, wire1356);
and AND3_473 (wire1359, n_63, n205, n273);
and AND3_474 (wire1360, n_62, n273, n86);
and AND3_475 (wire1361, n_61, n239, n273);
and AND3_476 (wire1362, n_60, n52, n273);
and AND3_477 (wire1363, n_59, n273, n35);
and AND3_478 (wire1364, n_58, n103, n273);
or OR2_479 (wire1368, wire1367, wire1366);
or OR2_480 (wire1372, wire1371, wire1370);
or OR2_481 (wire1376, wire1375, wire1374);
or OR2_482 (wire1380, wire1379, wire1378);
or OR2_483 (wire1384, wire1383, wire1382);
or OR2_484 (wire1388, wire1387, wire1386);
or OR2_485 (wire1392, wire1391, wire1390);
or OR2_486 (wire1396, wire1395, wire1394);
or OR2_487 (wire1400, wire1399, wire1398);
and AND3_488 (wire1401, n_47, n137, n273);
and AND3_489 (wire1402, n_46, n273, n69);
and AND3_490 (wire1403, n_45, n171, n273);
and AND3_491 (wire1404, n_44, n154, n273);
and AND3_492 (wire1405, n_43, n188, n273);
and AND3_493 (wire1406, n_42, n18, n273);
and AND3_494 (wire1407, n_41, n222, n273);
and AND3_495 (wire1408, n_40, n120, n273);
and AND2_496 (wire1412, wire1411, wire1409);
and AND2_497 (wire1416, wire1415, wire1413);
and AND2_498 (wire1420, wire1419, wire1417);
and AND2_499 (wire1424, wire1423, wire1421);
and AND2_500 (wire1428, wire1427, wire1425);
and AND2_501 (wire1432, wire1431, wire1429);
not NOT1_502 (n_711, wire1433);
not NOT1_503 (n_1290, wire1434);
not NOT1_504 (n_1075, wire1435);
not NOT1_505 (n_725, wire1436);
not NOT1_506 (n_447, wire1437);
not NOT1_507 (n_990, wire1438);
not NOT1_508 (n_168, wire1439);
not NOT1_509 (n_883, wire1440);
not NOT1_510 (n_731, wire1441);
not NOT1_511 (n_1026, wire1442);
not NOT1_512 (n_709, wire1443);
not NOT1_513 (n_994, wire1444);
not NOT1_514 (n_449, wire1445);
not NOT1_515 (n_1322, wire1446);
not NOT1_516 (n_1253, wire1447);
not NOT1_517 (n_1358, wire1448);
not NOT1_518 (n_740, wire1449);
not NOT1_519 (n_1341, wire1450);
not NOT1_520 (n_1114, wire1451);
not NOT1_521 (n_713, wire1452);
not NOT1_522 (n_368, wire1453);
not NOT1_523 (n_515, wire1454);
not NOT1_524 (n_1077, wire1455);
not NOT1_525 (n_1047, wire1456);
not NOT1_526 (n_1151, wire1457);
not NOT1_527 (n_1042, wire1458);
not NOT1_528 (n_267, wire1459);
not NOT1_529 (n_1404, wire1460);
not NOT1_530 (n_1107, wire1461);
not NOT1_531 (n_354, wire1462);
not NOT1_532 (n_1351, wire1463);
not NOT1_533 (n_1268, wire1464);
not NOT1_534 (n_360, wire1465);
not NOT1_535 (n_700, wire1466);
not NOT1_536 (n_548, wire1467);
not NOT1_537 (n_835, wire1468);
not NOT1_538 (n_461, wire1469);
not NOT1_539 (n_187, wire1470);
not NOT1_540 (n_455, wire1471);
not NOT1_541 (n_818, wire1472);
not NOT1_542 (n_191, wire1473);
not NOT1_543 (n_630, wire1474);
not NOT1_544 (n_362, wire1475);
not NOT1_545 (n_1144, wire1476);
not NOT1_546 (n_544, wire1477);
not NOT1_547 (n_808, wire1478);
not NOT1_548 (n_261, wire1479);
not NOT1_549 (n_1332, wire1480);
not NOT1_550 (n_562, wire1481);
not NOT1_551 (n_541, wire1482);
not NOT1_552 (n_257, wire1483);
not NOT1_553 (n_1336, wire1484);
not NOT1_554 (n_1424, wire1485);
not NOT1_555 (n_554, wire1486);
not NOT1_556 (n_166, wire1487);
not NOT1_557 (n_459, wire1488);
not NOT1_558 (n_350, wire1489);
not NOT1_559 (n_751, wire1490);
not NOT1_560 (n_1090, wire1491);
not NOT1_561 (n_79, wire1492);
not NOT1_562 (n_366, wire1493);
not NOT1_563 (n_633, wire1494);
not NOT1_564 (n_621, wire1495);
not NOT1_565 (n_856, wire1496);
not NOT1_566 (n_720, wire1497);
not NOT1_567 (n_443, wire1498);
not NOT1_568 (n545, wire1499);
and AND2_569 (wire1503, wire1502, wire1500);
and AND2_570 (wire1507, wire1506, wire1504);
not NOT1_571 (n_263, wire1508);
not NOT1_572 (n_1390, wire1509);
not NOT1_573 (n_531, wire1510);
not NOT1_574 (n_810, wire1511);
not NOT1_575 (n_164, wire1512);
not NOT1_576 (n_897, wire1513);
not NOT1_577 (n_981, wire1514);
not NOT1_578 (n_1155, wire1515);
not NOT1_579 (n_259, wire1516);
not NOT1_580 (n_643, wire1517);
not NOT1_581 (n_273, wire1518);
not NOT1_582 (n_1073, wire1519);
not NOT1_583 (n_985, wire1520);
not NOT1_584 (n_635, wire1521);
not NOT1_585 (n_265, wire1522);
not NOT1_586 (n_1003, wire1523);
not NOT1_587 (n_637, wire1524);
not NOT1_588 (n_457, wire1525);
not NOT1_589 (n_348, wire1526);
not NOT1_590 (n_812, wire1527);
not NOT1_591 (n_1096, wire1528);
not NOT1_592 (n_539, wire1529);
not NOT1_593 (n_624, wire1530);
not NOT1_594 (n_1385, wire1531);
not NOT1_595 (n_1081, wire1532);
not NOT1_596 (n_374, wire1533);
not NOT1_597 (n_1128, wire1534);
not NOT1_598 (n_799, wire1535);
not NOT1_599 (n_723, wire1536);
not NOT1_600 (n_1013, wire1537);
not NOT1_601 (n_1310, wire1538);
not NOT1_602 (n_826, wire1539);
not NOT1_603 (n_533, wire1540);
not NOT1_604 (n_734, wire1541);
not NOT1_605 (n_1255, wire1542);
not NOT1_606 (n_282, wire1543);
not NOT1_607 (n_1406, wire1544);
not NOT1_608 (n_1369, wire1545);
not NOT1_609 (n_189, wire1546);
not NOT1_610 (n_893, wire1547);
not NOT1_611 (n_886, wire1548);
not NOT1_612 (n_441, wire1549);
not NOT1_613 (n_278, wire1550);
not NOT1_614 (n_535, wire1551);
not NOT1_615 (n_284, wire1552);
not NOT1_616 (n_1348, wire1553);
not NOT1_617 (n_172, wire1554);
not NOT1_618 (n_453, wire1555);
not NOT1_619 (n_321, wire1556);
not NOT1_620 (n_352, wire1557);
not NOT1_621 (n_1021, wire1558);
not NOT1_622 (n_1338, wire1559);
not NOT1_623 (n_646, wire1560);
not NOT1_624 (n_177, wire1561);
not NOT1_625 (n_1283, wire1562);
not NOT1_626 (n_845, wire1563);
not NOT1_627 (n_626, wire1564);
not NOT1_628 (n_546, wire1565);
not NOT1_629 (n_356, wire1566);
not NOT1_630 (n_170, wire1567);
not NOT1_631 (n_901, wire1568);
not NOT1_632 (n_179, wire1569);
not NOT1_633 (n_1139, wire1570);
not NOT1_634 (n_801, wire1571);
not NOT1_635 (n_1432, wire1572);
not NOT1_636 (n_1300, wire1573);
not NOT1_637 (n_1439, wire1574);
not NOT1_638 (n_445, wire1575);
not NOT1_639 (n_656, wire1576);
not NOT1_640 (n_996, wire1577);
or OR2_641 (n_1524, wire1671, wire1670);
or OR2_642 (n_1525, wire1675, wire1674);
not NOT1_643 (wire1758, n_34);
not NOT1_644 (wire1121, n_996);
and AND2_645 (wire1301, n_79, n_100);
not NOT1_646 (n_80, wire1313);
or OR2_647 (wire1314, n_79, n_100);
not NOT1_648 (n_78, wire1318);
not NOT1_649 (n_76, wire1322);
not NOT1_650 (n_75, wire1326);
not NOT1_651 (n_74, wire1330);
not NOT1_652 (n_72, wire1334);
not NOT1_653 (n_71, wire1338);
not NOT1_654 (n_70, wire1342);
not NOT1_655 (n_69, wire1346);
not NOT1_656 (n_68, wire1350);
not NOT1_657 (n_66, wire1354);
not NOT1_658 (n_65, wire1358);
not NOT1_659 (n_98, wire1359);
not NOT1_660 (n_82, wire1360);
not NOT1_661 (n_86, wire1361);
not NOT1_662 (n_83, wire1362);
not NOT1_663 (n_91, wire1363);
not NOT1_664 (n_92, wire1364);
not NOT1_665 (n_57, wire1368);
not NOT1_666 (n_56, wire1372);
not NOT1_667 (n_55, wire1376);
not NOT1_668 (n_54, wire1380);
not NOT1_669 (n_53, wire1384);
not NOT1_670 (n_52, wire1388);
not NOT1_671 (n_51, wire1392);
not NOT1_672 (n_50, wire1396);
not NOT1_673 (n_49, wire1400);
not NOT1_674 (n_97, wire1401);
not NOT1_675 (n_85, wire1402);
not NOT1_676 (n_95, wire1403);
not NOT1_677 (n_84, wire1404);
not NOT1_678 (n_81, wire1405);
not NOT1_679 (n_94, wire1406);
not NOT1_680 (n_96, wire1407);
not NOT1_681 (n_93, wire1408);
not NOT1_682 (n_39, wire1412);
not NOT1_683 (n_38, wire1416);
not NOT1_684 (n_37, wire1420);
not NOT1_685 (n_36, wire1424);
not NOT1_686 (n_33, wire1428);
not NOT1_687 (n_32, wire1432);
not NOT1_688 (n_7, wire1503);
not NOT1_689 (n_6, wire1507);
or OR2_690 (wire1122, wire1121, n_888);
and AND2_691 (wire1267, n_92, n_58);
and AND2_692 (wire1269, n_94, n_42);
and AND2_693 (wire1271, n_83, n_60);
and AND2_694 (wire1273, n_98, n_63);
and AND2_695 (wire1275, n_97, n_47);
and AND2_696 (wire1277, n_91, n_59);
and AND2_697 (wire1278, n_81, n_43);
and AND2_698 (wire1280, n_93, n_40);
and AND2_699 (wire1281, n_95, n_45);
and AND4_700 (wire1283, n_80, n_77, n_23, n_27);
and AND2_701 (wire1284, n_85, n_46);
and AND2_702 (wire1287, n_84, n_44);
and AND2_703 (wire1289, n_96, n_41);
and AND2_704 (wire1291, n_86, n_61);
and AND2_705 (wire1293, n_82, n_62);
and AND4_706 (wire1295, n_1524, n_68, n_65, n_6);
and AND4_707 (wire1296, n_53, n_74, n_78, n_37);
and AND4_708 (wire1297, n_72, n_1525, n_69, n_7);
and AND4_709 (wire1298, n_51, n_70, n_32, n_33);
and AND4_710 (wire1299, n_54, n_52, n_76, n_39);
and AND4_711 (wire1300, n_57, n_50, n_36, n_38);
and AND3_712 (n_122, n_98, n205, n273);
and AND3_713 (n_129, n_97, n137, n273);
and AND3_714 (n_114, n_96, n222, n273);
and AND3_715 (n_131, n_95, n171, n273);
and AND3_716 (wire1302, n_94, n18, n273);
and AND3_717 (n_135, n_93, n120, n273);
and AND3_718 (wire1303, n_92, n103, n273);
and AND3_719 (n_141, n_91, n273, n35);
and AND2_720 (wire1307, wire1306, n_71);
and AND2_721 (wire1311, wire1310, n_49);
and AND3_722 (n_113, n_86, n239, n273);
and AND3_723 (n_133, n_85, n69, n273);
and AND3_724 (n_139, n_84, n154, n273);
and AND3_725 (wire1312, n_83, n52, n273);
and AND3_726 (n_145, n_82, n86, n273);
and AND3_727 (n_137, n_81, n188, n273);
not NOT1_728 (n_99, wire1314);
or OR2_729 (wire1123, wire1122, n_1153);
or OR2_730 (wire1274, wire1273, n_122);
or OR2_731 (wire1276, wire1275, n_129);
or OR2_732 (n_117, wire1277, n_141);
or OR2_733 (wire1279, wire1278, n_137);
or OR2_734 (n_121, wire1280, n_135);
or OR2_735 (wire1282, wire1281, n_131);
not NOT1_736 (n_110, wire1283);
or OR2_737 (n_119, wire1284, n_133);
or OR2_738 (wire1285, n_100, n_99);
or OR2_739 (wire1288, wire1287, n_139);
or OR2_740 (wire1290, wire1289, n_114);
or OR2_741 (wire1292, wire1291, n_113);
or OR2_742 (wire1294, wire1293, n_145);
not NOT1_743 (n_109, wire1295);
not NOT1_744 (n_108, wire1296);
not NOT1_745 (n_106, wire1297);
not NOT1_746 (n_105, wire1298);
not NOT1_747 (n_103, wire1299);
not NOT1_748 (n_102, wire1300);
or OR2_749 (n_112, wire1301, n_99);
not NOT1_750 (n_116, wire1302);
not NOT1_751 (n_120, wire1303);
not NOT1_752 (n_90, wire1307);
not NOT1_753 (n_88, wire1311);
not NOT1_754 (n_118, wire1312);
or OR2_755 (wire1235, n_117, n_116);
or OR2_756 (wire1237, n_121, n_120);
or OR2_757 (wire1245, n_119, n_118);
and AND2_758 (wire1247, n_113, n_112);
or OR4_759 (wire1249, n_110, n_67, n205, n137);
or OR4_760 (wire1258, n_106, n_90, n_75, n_66);
or OR4_761 (wire1259, n_102, n_88, n_56, n_55);
or OR4_762 (wire1260, n_108, n_109, n_103, n_105);
and AND2_763 (wire1262, n_121, n_120);
and AND2_764 (wire1263, n_119, n_118);
and AND2_765 (wire1264, n_117, n_116);
or OR2_766 (wire1266, n_113, n_112);
not NOT1_767 (n_138, wire1274);
not NOT1_768 (n_136, wire1276);
not NOT1_769 (n_132, wire1279);
not NOT1_770 (n_140, wire1282);
and AND2_771 (wire1286, wire1285, n290);
not NOT1_772 (n_130, wire1288);
not NOT1_773 (n_123, wire1290);
not NOT1_774 (n_115, wire1292);
not NOT1_775 (n_134, wire1294);
not NOT1_776 (n_107, n_120);
not NOT1_777 (n_104, n_116);
not NOT1_778 (n_101, n_118);
and AND2_779 (wire1233, n_123, n_122);
and AND2_780 (wire1234, n_130, n_129);
and AND2_781 (wire1236, n_138, n_137);
and AND2_782 (wire1238, n_134, n_133);
and AND2_783 (wire1239, n_115, n_114);
and AND2_784 (wire1240, n_132, n_131);
and AND2_785 (wire1241, n_140, n_139);
and AND2_786 (wire1244, n_136, n_135);
not NOT1_787 (n_143, wire1249);
or OR2_788 (wire1251, n_140, n_139);
or OR2_789 (wire1252, n_138, n_137);
or OR2_790 (wire1253, n_136, n_135);
or OR2_791 (wire1254, n_134, n_133);
or OR2_792 (wire1255, n_132, n_131);
or OR2_793 (wire1256, n_130, n_129);
not NOT1_794 (n_126, wire1258);
not NOT1_795 (n_125, wire1259);
not NOT1_796 (n_124, wire1260);
or OR2_797 (wire1261, n_123, n_122);
not NOT1_798 (n_155, wire1262);
not NOT1_799 (n_147, wire1263);
not NOT1_800 (n_157, wire1264);
or OR2_801 (wire1265, n_115, n_114);
not NOT1_802 (n_144, wire1266);
or OR2_803 (wire1268, wire1267, n_107);
or OR2_804 (wire1270, wire1269, n_104);
or OR2_805 (wire1272, wire1271, n_101);
and AND2_806 (n_128, wire1286, n256);
and AND2_807 (wire1035, n_124, n_125);
and AND4_808 (wire1224, n_143, n_73, n358, n341);
and AND2_809 (n_184, wire1235, n_157);
and AND2_810 (n_186, wire1237, n_155);
or OR2_811 (wire1242, n_128, n_127);
and AND2_812 (n_182, wire1245, n_147);
or OR2_813 (wire1248, wire1247, n_144);
not NOT1_814 (n_149, wire1251);
not NOT1_815 (n_156, wire1252);
not NOT1_816 (n_148, wire1253);
not NOT1_817 (n_154, wire1254);
not NOT1_818 (n_150, wire1255);
not NOT1_819 (n_158, wire1256);
and AND2_820 (wire1257, n_128, n_127);
not NOT1_821 (n_159, wire1261);
not NOT1_822 (n_151, wire1265);
not NOT1_823 (n_146, wire1268);
not NOT1_824 (n1581, wire1270);
not NOT1_825 (n_142, wire1272);
and AND2_826 (wire1036, wire1035, n_126);
or OR2_827 (wire1185, n_184, n_183);
or OR2_828 (wire1192, n_182, n_181);
or OR2_829 (wire1206, n_186, n_185);
and AND2_830 (wire1219, n_186, n_185);
and AND2_831 (wire1220, n_184, n_183);
and AND2_832 (wire1221, n_182, n_181);
not NOT1_833 (n_174, wire1224);
and AND2_834 (wire1230, n_142, n_141);
and AND2_835 (wire1232, n_146, n_145);
or OR2_836 (n_167, wire1233, n_159);
or OR2_837 (n_171, wire1234, n_158);
or OR2_838 (n_180, wire1236, n_156);
or OR2_839 (n_169, wire1238, n_154);
or OR2_840 (n_178, wire1239, n_151);
or OR2_841 (n_165, wire1240, n_150);
or OR2_842 (n_173, wire1241, n_149);
or OR2_843 (n_188, wire1244, n_148);
or OR2_844 (wire1246, n_146, n_145);
not NOT1_845 (n_162, wire1248);
or OR2_846 (wire1250, n_142, n_141);
not NOT1_847 (n_152, wire1257);
or OR4_848 (wire1176, n_174, n307, n222, n154);
and AND2_849 (wire1178, n_152, n290);
and AND2_850 (wire1187, n_169, n_168);
and AND2_851 (wire1189, n_178, n_177);
and AND2_852 (wire1190, n_165, n_164);
and AND2_853 (wire1191, n_171, n_170);
and AND2_854 (wire1195, n_173, n_172);
and AND2_855 (wire1208, n_188, n_187);
and AND2_856 (wire1210, n_180, n_179);
and AND2_857 (wire1211, n_167, n_166);
or OR2_858 (wire1216, n_162, n_161);
or OR2_859 (wire1218, n_188, n_187);
not NOT1_860 (n_196, wire1219);
not NOT1_861 (n_202, wire1220);
not NOT1_862 (n_203, wire1221);
or OR2_863 (wire1222, n_180, n_179);
or OR2_864 (wire1223, n_178, n_177);
or OR2_865 (wire1225, n_173, n_172);
or OR2_866 (wire1226, n_171, n_170);
or OR2_867 (wire1227, n_169, n_168);
or OR2_868 (wire1228, n_167, n_166);
or OR2_869 (wire1229, n_165, n_164);
and AND2_870 (wire1231, n_162, n_161);
and AND2_871 (n_153, n_152, n290);
and AND2_872 (wire1243, wire1242, n_152);
not NOT1_873 (n_160, wire1246);
not NOT1_874 (n_163, wire1250);
not NOT1_875 (n_208, wire1176);
and AND2_876 (wire1179, wire1178, n307);
and AND2_877 (wire1186, wire1185, n_202);
and AND2_878 (wire1193, wire1192, n_203);
and AND2_879 (wire1196, n_203, n_147);
and AND2_880 (wire1197, n_202, n_157);
and AND2_881 (wire1205, n_196, n_155);
and AND2_882 (wire1207, wire1206, n_196);
or OR2_883 (wire1214, n_153, n307);
not NOT1_884 (n_195, wire1218);
not NOT1_885 (n_194, wire1222);
not NOT1_886 (n_198, wire1223);
not NOT1_887 (n_201, wire1225);
not NOT1_888 (n_199, wire1226);
not NOT1_889 (n_200, wire1227);
not NOT1_890 (n_193, wire1228);
not NOT1_891 (n_197, wire1229);
or OR2_892 (n_190, wire1230, n_163);
not NOT1_893 (n_175, wire1231);
or OR2_894 (n_192, wire1232, n_160);
not NOT1_895 (n_209, wire1243);
and AND4_896 (wire1149, n_208, n_89, n_15, n392);
and AND2_897 (wire1177, n_192, n_191);
and AND2_898 (wire1183, n_190, n_189);
not NOT1_899 (n1901, wire1186);
or OR2_900 (wire1188, wire1187, n_200);
or OR2_901 (n_216, wire1189, n_198);
or OR2_902 (n_222, wire1190, n_197);
or OR2_903 (n_226, wire1191, n_199);
not NOT1_904 (n_232, wire1193);
or OR2_905 (wire1194, n_193, n_159);
or OR2_906 (n_220, wire1195, n_201);
not NOT1_907 (n_223, wire1196);
not NOT1_908 (n_236, wire1197);
or OR2_909 (wire1198, n_201, n_149);
or OR2_910 (wire1199, n_200, n_154);
or OR2_911 (wire1200, n_199, n_158);
or OR2_912 (wire1201, n_198, n_151);
or OR2_913 (wire1202, n_194, n_156);
or OR2_914 (wire1203, n_195, n_148);
or OR2_915 (wire1204, n_197, n_150);
not NOT1_916 (n_227, wire1205);
not NOT1_917 (n_238, wire1207);
or OR2_918 (wire1209, wire1208, n_195);
or OR2_919 (n_214, wire1210, n_194);
or OR2_920 (n_218, wire1211, n_193);
or OR2_921 (wire1212, n_192, n_191);
or OR2_922 (wire1213, n_190, n_189);
and AND2_923 (wire1215, wire1214, n256);
and AND2_924 (wire1217, wire1216, n_175);
not NOT1_925 (wire1756, n_175);
not NOT1_926 (n_249, wire1149);
not NOT1_927 (n_224, wire1188);
not NOT1_928 (n_215, wire1194);
not NOT1_929 (n_221, wire1198);
not NOT1_930 (n_229, wire1199);
not NOT1_931 (n_219, wire1200);
not NOT1_932 (n_212, wire1201);
not NOT1_933 (n_217, wire1202);
not NOT1_934 (n_225, wire1203);
not NOT1_935 (n_213, wire1204);
not NOT1_936 (n_228, wire1209);
not NOT1_937 (n_206, wire1212);
not NOT1_938 (n_205, wire1213);
not NOT1_939 (n_207, wire1215);
not NOT1_940 (n_211, wire1217);
or OR2_941 (wire1757, wire1756, n_144);
or OR2_942 (wire1124, wire1123, n_249);
and AND2_943 (wire1150, n_214, n_213);
and AND2_944 (wire1151, n_218, n_217);
and AND2_945 (wire1152, n_212, n_211);
or OR2_946 (wire1153, n_228, n_227);
or OR2_947 (wire1154, n_224, n_223);
and AND2_948 (wire1155, n_220, n_219);
and AND2_949 (wire1156, n_216, n_215);
and AND2_950 (wire1157, n_226, n_225);
and AND2_951 (wire1158, n_222, n_221);
and AND2_952 (wire1166, n_228, n_227);
or OR2_953 (wire1167, n_226, n_225);
and AND2_954 (wire1168, n_224, n_223);
or OR2_955 (wire1169, n_222, n_221);
or OR2_956 (wire1170, n_220, n_219);
or OR2_957 (wire1171, n_218, n_217);
or OR2_958 (wire1172, n_216, n_215);
or OR2_959 (wire1173, n_214, n_213);
or OR2_960 (wire1174, n_212, n_211);
or OR2_961 (n_230, wire1177, n_206);
or OR2_962 (wire1180, wire1179, n_207);
or OR2_963 (wire1181, n_206, n_160);
or OR2_964 (wire1182, n_205, n_163);
or OR2_965 (wire1184, wire1183, n_205);
not NOT1_966 (n_1566, wire1757);
not NOT1_967 (n_286, wire1124);
and AND2_968 (wire1142, n_230, n_229);
and AND2_969 (wire1159, n_1566, n_209);
or OR2_970 (wire1165, n_230, n_229);
not NOT1_971 (n_245, wire1166);
not NOT1_972 (n_241, wire1167);
not NOT1_973 (n_244, wire1168);
not NOT1_974 (n_240, wire1169);
not NOT1_975 (n_243, wire1170);
not NOT1_976 (n_247, wire1171);
not NOT1_977 (n_242, wire1172);
not NOT1_978 (n_248, wire1173);
not NOT1_979 (n_246, wire1174);
or OR2_980 (wire1175, n_1566, n_209);
not NOT1_981 (n_234, wire1180);
not NOT1_982 (n_237, wire1181);
not NOT1_983 (n_231, wire1182);
not NOT1_984 (n_235, wire1184);
and AND4_985 (wire1077, n_286, n_18, n_87, n103);
and AND2_986 (wire1141, n_232, n_231);
or OR2_987 (wire1145, n_236, n_235);
or OR2_988 (wire1146, n_234, n_233);
and AND2_989 (wire1148, n_238, n_237);
or OR2_990 (n_274, wire1150, n_248);
or OR2_991 (n_264, wire1151, n_247);
or OR2_992 (n_262, wire1152, n_246);
and AND2_993 (n_272, wire1153, n_245);
and AND2_994 (n_270, wire1154, n_244);
or OR2_995 (n_260, wire1155, n_243);
or OR2_996 (n_266, wire1156, n_242);
or OR2_997 (n_268, wire1157, n_241);
or OR2_998 (n_258, wire1158, n_240);
or OR2_999 (wire1161, n_238, n_237);
and AND2_1000 (wire1162, n_236, n_235);
and AND2_1001 (wire1163, n_234, n_233);
or OR2_1002 (wire1164, n_232, n_231);
not NOT1_1003 (n_253, wire1165);
not NOT1_1004 (n_239, wire1175);
not NOT1_1005 (n_318, wire1077);
or OR2_1006 (wire1107, n_272, n_271);
or OR2_1007 (wire1109, n_270, n_269);
and AND2_1008 (wire1111, n_258, n_257);
and AND2_1009 (wire1112, n_262, n_261);
and AND2_1010 (wire1113, n_274, n_273);
and AND2_1011 (wire1114, n_268, n_267);
and AND2_1012 (wire1116, n_264, n_263);
and AND2_1013 (wire1117, n_266, n_265);
and AND2_1014 (wire1118, n_260, n_259);
or OR2_1015 (wire1131, n_274, n_273);
and AND2_1016 (wire1132, n_272, n_271);
and AND2_1017 (wire1133, n_270, n_269);
or OR2_1018 (wire1134, n_268, n_267);
or OR2_1019 (wire1135, n_266, n_265);
or OR2_1020 (wire1136, n_264, n_263);
or OR2_1021 (wire1137, n_262, n_261);
or OR2_1022 (wire1138, n_260, n_259);
or OR2_1023 (wire1139, n_258, n_257);
or OR2_1024 (n_283, wire1142, n_253);
or OR2_1025 (wire1160, wire1159, n_239);
not NOT1_1026 (n_250, wire1161);
not NOT1_1027 (n_252, wire1162);
not NOT1_1028 (n_251, wire1163);
not NOT1_1029 (n_254, wire1164);
or OR4_1030 (wire1054, n_318, n477, n426, n409);
and AND2_1031 (wire1093, n_283, n_282);
or OR2_1032 (wire1126, n_283, n_282);
not NOT1_1033 (n_291, wire1131);
not NOT1_1034 (n_295, wire1132);
not NOT1_1035 (n_294, wire1133);
not NOT1_1036 (n_290, wire1134);
not NOT1_1037 (n_288, wire1135);
not NOT1_1038 (n_289, wire1136);
not NOT1_1039 (n_292, wire1137);
not NOT1_1040 (n_287, wire1138);
not NOT1_1041 (n_293, wire1139);
or OR2_1042 (n_279, wire1141, n_254);
not NOT1_1043 (wire1143, n_251);
and AND2_1044 (n_277, wire1145, n_252);
and AND2_1045 (wire1147, wire1146, n_251);
or OR2_1046 (n_285, wire1148, n_250);
not NOT1_1047 (n_256, wire1160);
not NOT1_1048 (n_373, wire1054);
and AND2_1049 (wire1090, n_285, n_284);
or OR2_1050 (wire1091, n_277, n_276);
and AND2_1051 (wire1095, n_279, n_278);
and AND2_1052 (wire1098, n_294, n_244);
or OR2_1053 (wire1099, n_288, n_242);
or OR2_1054 (wire1100, n_293, n_240);
or OR2_1055 (wire1101, n_292, n_246);
or OR2_1056 (wire1102, n_291, n_248);
or OR2_1057 (wire1103, n_289, n_247);
or OR2_1058 (wire1104, n_290, n_241);
or OR2_1059 (wire1105, n_287, n_243);
and AND2_1060 (wire1106, n_295, n_245);
and AND2_1061 (wire1108, wire1107, n_295);
and AND2_1062 (wire1110, wire1109, n_294);
or OR2_1063 (n_309, wire1111, n_293);
or OR2_1064 (n_312, wire1112, n_292);
or OR2_1065 (n_303, wire1113, n_291);
or OR2_1066 (wire1115, wire1114, n_290);
or OR2_1067 (n_311, wire1116, n_289);
or OR2_1068 (n_307, wire1117, n_288);
or OR2_1069 (n_305, wire1118, n_287);
or OR2_1070 (wire1119, n_256, n_255);
or OR2_1071 (wire1125, n_285, n_284);
not NOT1_1072 (n_298, wire1126);
or OR2_1073 (wire1127, n_279, n_278);
and AND2_1074 (wire1128, n_277, n_276);
and AND2_1075 (wire1140, n_256, n_255);
or OR2_1076 (wire1144, wire1143, n_207);
not NOT1_1077 (n_319, wire1147);
or OR2_1078 (wire1037, wire1036, n_373);
or OR2_1079 (wire1086, n_298, n_253);
or OR2_1080 (wire1094, wire1093, n_298);
not NOT1_1081 (n_327, wire1098);
not NOT1_1082 (n_313, wire1099);
not NOT1_1083 (n_302, wire1100);
not NOT1_1084 (n_317, wire1101);
not NOT1_1085 (n_310, wire1102);
not NOT1_1086 (n_306, wire1103);
not NOT1_1087 (n_304, wire1104);
not NOT1_1088 (n_308, wire1105);
not NOT1_1089 (n_314, wire1106);
not NOT1_1090 (n_330, wire1108);
not NOT1_1091 (n_324, wire1110);
not NOT1_1092 (n_315, wire1115);
not NOT1_1093 (n_301, wire1125);
not NOT1_1094 (n_297, wire1127);
not NOT1_1095 (n_299, wire1128);
not NOT1_1096 (n_280, wire1140);
not NOT1_1097 (n_275, wire1144);
not NOT1_1098 (n_1412, wire1037);
and AND2_1099 (wire1062, n_303, n_302);
and AND2_1100 (wire1063, n_311, n_310);
and AND2_1101 (wire1064, n_313, n_312);
and AND2_1102 (wire1066, n_307, n_306);
and AND2_1103 (wire1067, n_309, n_308);
and AND2_1104 (wire1068, n_305, n_304);
or OR2_1105 (wire1069, n_315, n_314);
and AND2_1106 (wire1079, n_315, n_314);
or OR2_1107 (wire1080, n_313, n_312);
or OR2_1108 (wire1081, n_311, n_310);
or OR2_1109 (wire1082, n_309, n_308);
or OR2_1110 (wire1083, n_307, n_306);
or OR2_1111 (wire1084, n_305, n_304);
or OR2_1112 (wire1085, n_303, n_302);
not NOT1_1113 (n_325, wire1086);
or OR2_1114 (wire1087, n_301, n_250);
and AND2_1115 (wire1088, n_299, n_252);
or OR2_1116 (wire1089, n_297, n_254);
or OR2_1117 (n_326, wire1090, n_301);
and AND2_1118 (wire1092, wire1091, n_299);
not NOT1_1119 (n_328, wire1094);
or OR2_1120 (wire1096, wire1095, n_297);
and AND2_1121 (wire1097, n_275, n324);
and AND2_1122 (wire1120, wire1119, n_280);
or OR2_1123 (wire1130, wire1129, n_275);
not NOT1_1124 (wire1754, n_280);
or OR2_1125 (wire1055, n_328, n_327);
and AND2_1126 (wire1058, n_326, n_325);
and AND2_1127 (wire1072, n_328, n_327);
or OR2_1128 (wire1073, n_326, n_325);
not NOT1_1129 (n_333, wire1079);
not NOT1_1130 (n_338, wire1080);
not NOT1_1131 (n_339, wire1081);
not NOT1_1132 (n_335, wire1082);
not NOT1_1133 (n_336, wire1083);
not NOT1_1134 (n_334, wire1084);
not NOT1_1135 (n_340, wire1085);
not NOT1_1136 (n_329, wire1087);
not NOT1_1137 (n_332, wire1088);
not NOT1_1138 (n_323, wire1089);
not NOT1_1139 (n2223, wire1092);
not NOT1_1140 (n_331, wire1096);
not NOT1_1141 (n_316, wire1120);
not NOT1_1142 (n_296, wire1130);
or OR2_1143 (wire1755, wire1754, n_239);
and AND2_1144 (wire1052, n_330, n_329);
or OR2_1145 (wire1057, n_332, n_331);
and AND2_1146 (wire1059, n_324, n_323);
or OR2_1147 (n_349, wire1062, n_340);
or OR2_1148 (n_353, wire1063, n_339);
or OR2_1149 (n_363, wire1064, n_338);
and AND2_1150 (wire1065, n_317, n_316);
or OR2_1151 (n_351, wire1066, n_336);
or OR2_1152 (n_361, wire1067, n_335);
or OR2_1153 (n_357, wire1068, n_334);
and AND2_1154 (n_359, wire1069, n_333);
and AND2_1155 (wire1070, n_332, n_331);
or OR2_1156 (wire1071, n_330, n_329);
not NOT1_1157 (n_346, wire1072);
not NOT1_1158 (n_343, wire1073);
or OR2_1159 (wire1074, n_324, n_323);
or OR2_1160 (wire1078, n_317, n_316);
or OR2_1161 (n_322, wire1097, n_296);
not NOT1_1162 (n_1565, wire1755);
and AND2_1163 (wire1023, n_351, n_350);
and AND2_1164 (wire1025, n_361, n_360);
and AND2_1165 (wire1026, n_353, n_352);
and AND2_1166 (wire1027, n_349, n_348);
and AND2_1167 (wire1028, n_357, n_356);
or OR2_1168 (wire1030, n_359, n_358);
and AND2_1169 (wire1032, n_363, n_362);
or OR2_1170 (wire1044, n_363, n_362);
or OR2_1171 (wire1045, n_361, n_360);
and AND2_1172 (wire1046, n_359, n_358);
or OR2_1173 (wire1047, n_357, n_356);
or OR2_1174 (wire1049, n_353, n_352);
or OR2_1175 (wire1050, n_351, n_350);
or OR2_1176 (wire1051, n_349, n_348);
and AND2_1177 (n_372, wire1055, n_346);
and AND2_1178 (wire1056, n_322, n_321);
or OR2_1179 (n_369, wire1058, n_343);
and AND2_1180 (wire1060, n_1565, n_319);
not NOT1_1181 (n_344, wire1070);
not NOT1_1182 (n_347, wire1071);
not NOT1_1183 (n_342, wire1074);
or OR2_1184 (wire1075, n_322, n_321);
or OR2_1185 (wire1076, n_1565, n_319);
not NOT1_1186 (n_337, wire1078);
or OR2_1187 (wire1004, n_372, n_371);
and AND2_1188 (wire1006, n_369, n_368);
and AND2_1189 (wire1038, n_372, n_371);
or OR2_1190 (wire1041, n_369, n_368);
not NOT1_1191 (n_378, wire1044);
not NOT1_1192 (n_383, wire1045);
not NOT1_1193 (n_379, wire1046);
not NOT1_1194 (n_380, wire1047);
not NOT1_1195 (n_382, wire1049);
not NOT1_1196 (n_385, wire1050);
not NOT1_1197 (n_381, wire1051);
or OR2_1198 (n_375, wire1052, n_347);
and AND2_1199 (n_377, wire1057, n_344);
or OR2_1200 (n_367, wire1059, n_342);
or OR2_1201 (n_355, wire1065, n_337);
not NOT1_1202 (n_345, wire1075);
not NOT1_1203 (n_341, wire1076);
or OR2_1204 (wire997, n_377, n_376);
and AND2_1205 (wire1008, n_375, n_374);
and AND2_1206 (wire1009, n_367, n_366);
or OR2_1207 (wire1016, n_385, n_336);
or OR2_1208 (wire1017, n_383, n_335);
or OR2_1209 (wire1018, n_378, n_338);
and AND2_1210 (wire1019, n_379, n_333);
or OR2_1211 (wire1020, n_381, n_340);
or OR2_1212 (wire1021, n_382, n_339);
or OR2_1213 (wire1022, n_380, n_334);
or OR2_1214 (n_396, wire1023, n_385);
and AND2_1215 (wire1024, n_355, n_354);
or OR2_1216 (n_406, wire1025, n_383);
or OR2_1217 (n_398, wire1026, n_382);
or OR2_1218 (n_400, wire1027, n_381);
or OR2_1219 (wire1029, wire1028, n_380);
and AND2_1220 (wire1031, wire1030, n_379);
or OR2_1221 (n_408, wire1032, n_378);
and AND2_1222 (wire1033, n_377, n_376);
or OR2_1223 (wire1034, n_375, n_374);
not NOT1_1224 (n_392, wire1038);
not NOT1_1225 (n_391, wire1041);
or OR2_1226 (wire1042, n_367, n_366);
or OR2_1227 (wire1048, n_355, n_354);
or OR2_1228 (wire1053, n_345, n_296);
or OR2_1229 (n_423, wire1056, n_345);
or OR2_1230 (wire1061, wire1060, n_341);
and AND2_1231 (wire1000, n_392, n_346);
or OR2_1232 (wire1003, n_391, n_343);
and AND2_1233 (wire1005, wire1004, n_392);
or OR2_1234 (wire1007, wire1006, n_391);
not NOT1_1235 (n_407, wire1016);
not NOT1_1236 (n_399, wire1017);
not NOT1_1237 (n_402, wire1018);
not NOT1_1238 (n_403, wire1019);
not NOT1_1239 (n_397, wire1020);
not NOT1_1240 (n_395, wire1021);
not NOT1_1241 (n_405, wire1022);
not NOT1_1242 (n_404, wire1029);
not NOT1_1243 (n_422, wire1031);
not NOT1_1244 (n_393, wire1033);
not NOT1_1245 (n_390, wire1034);
not NOT1_1246 (n_389, wire1042);
not NOT1_1247 (n_384, wire1048);
not NOT1_1248 (n_370, wire1053);
not NOT1_1249 (n_365, wire1061);
and AND2_1250 (wire975, n_400, n_399);
and AND2_1251 (wire976, n_408, n_407);
and AND2_1252 (wire977, n_398, n_397);
and AND2_1253 (wire979, n_396, n_395);
or OR2_1254 (wire980, n_404, n_403);
and AND2_1255 (wire981, n_406, n_405);
or OR2_1256 (wire990, n_408, n_407);
or OR2_1257 (wire991, n_406, n_405);
and AND2_1258 (wire992, n_404, n_403);
or OR2_1259 (wire994, n_400, n_399);
or OR2_1260 (wire995, n_398, n_397);
or OR2_1261 (wire996, n_396, n_395);
and AND2_1262 (wire998, wire997, n_393);
or OR2_1263 (wire999, n_390, n_347);
not NOT1_1264 (n_419, wire1000);
and AND2_1265 (wire1001, n_393, n_344);
or OR2_1266 (wire1002, n_389, n_342);
not NOT1_1267 (n_409, wire1003);
not NOT1_1268 (n_416, wire1005);
not NOT1_1269 (n_420, wire1007);
or OR2_1270 (n_410, wire1008, n_390);
or OR2_1271 (wire1010, wire1009, n_389);
and AND2_1272 (wire1011, n_370, n341);
or OR2_1273 (wire1013, n_365, n_364);
or OR2_1274 (wire1015, n_384, n_337);
or OR2_1275 (n_401, wire1024, n_384);
or OR2_1276 (wire1040, wire1039, n_370);
and AND2_1277 (wire1043, n_365, n_364);
and AND2_1278 (wire971, n_410, n_409);
or OR2_1279 (wire973, n_420, n_419);
and AND2_1280 (wire978, n_402, n_401);
and AND2_1281 (wire984, n_420, n_419);
or OR2_1282 (wire989, n_410, n_409);
not NOT1_1283 (n_432, wire990);
not NOT1_1284 (n_425, wire991);
not NOT1_1285 (n_426, wire992);
or OR2_1286 (wire993, n_402, n_401);
not NOT1_1287 (n_433, wire994);
not NOT1_1288 (n_431, wire995);
not NOT1_1289 (n_427, wire996);
not NOT1_1290 (n2548, wire998);
not NOT1_1291 (n_421, wire999);
not NOT1_1292 (n_418, wire1001);
not NOT1_1293 (n_415, wire1002);
not NOT1_1294 (n_417, wire1010);
not NOT1_1295 (n_414, wire1015);
not NOT1_1296 (n_388, wire1040);
not NOT1_1297 (n_386, wire1043);
and AND2_1298 (wire967, n_416, n_415);
or OR2_1299 (wire970, n_418, n_417);
and AND2_1300 (wire972, n_422, n_421);
or OR2_1301 (n_454, wire975, n_433);
or OR2_1302 (n_446, wire976, n_432);
or OR2_1303 (n_444, wire977, n_431);
or OR2_1304 (n_450, wire979, n_427);
and AND2_1305 (n_452, wire980, n_426);
or OR2_1306 (n_442, wire981, n_425);
or OR2_1307 (wire983, n_422, n_421);
not NOT1_1308 (n_435, wire984);
and AND2_1309 (wire985, n_418, n_417);
or OR2_1310 (wire986, n_416, n_415);
not NOT1_1311 (n_437, wire989);
not NOT1_1312 (n_430, wire993);
or OR2_1313 (wire1012, wire1011, n_388);
and AND2_1314 (wire1014, wire1013, n_386);
not NOT1_1315 (wire1752, n_386);
or OR2_1316 (wire940, n_452, n_451);
and AND2_1317 (wire942, n_444, n_443);
and AND2_1318 (wire943, n_446, n_445);
and AND2_1319 (wire944, n_454, n_453);
and AND2_1320 (wire946, n_442, n_441);
and AND2_1321 (wire948, n_450, n_449);
or OR2_1322 (wire958, n_454, n_453);
and AND2_1323 (wire959, n_452, n_451);
or OR2_1324 (wire960, n_450, n_449);
or OR2_1325 (wire962, n_446, n_445);
or OR2_1326 (wire963, n_444, n_443);
or OR2_1327 (wire964, n_442, n_441);
or OR2_1328 (n_460, wire971, n_437);
and AND2_1329 (n_464, wire973, n_435);
or OR2_1330 (n_448, wire978, n_430);
not NOT1_1331 (n_436, wire983);
not NOT1_1332 (n_438, wire985);
not NOT1_1333 (n_439, wire986);
not NOT1_1334 (n_412, wire1012);
not NOT1_1335 (n_413, wire1014);
or OR2_1336 (wire1753, wire1752, n_341);
and AND2_1337 (wire927, n_460, n_459);
or OR2_1338 (wire931, n_464, n_463);
and AND2_1339 (wire945, n_448, n_447);
and AND2_1340 (wire953, n_464, n_463);
or OR2_1341 (wire955, n_460, n_459);
not NOT1_1342 (n_473, wire958);
not NOT1_1343 (n_476, wire959);
not NOT1_1344 (n_470, wire960);
or OR2_1345 (wire961, n_448, n_447);
not NOT1_1346 (n_474, wire962);
not NOT1_1347 (n_475, wire963);
not NOT1_1348 (n_471, wire964);
or OR2_1349 (n_458, wire967, n_439);
or OR2_1350 (wire968, n_412, n_411);
and AND2_1351 (n_466, wire970, n_438);
or OR2_1352 (n_462, wire972, n_436);
and AND2_1353 (wire974, n_414, n_413);
or OR2_1354 (wire987, n_414, n_413);
and AND2_1355 (wire988, n_412, n_411);
not NOT1_1356 (n_1564, wire1753);
or OR2_1357 (wire923, n_466, n_465);
and AND2_1358 (wire925, n_458, n_457);
and AND2_1359 (wire930, n_462, n_461);
or OR2_1360 (wire933, n_473, n_433);
or OR2_1361 (wire934, n_470, n_427);
or OR2_1362 (wire935, n_471, n_425);
or OR2_1363 (wire936, n_474, n_432);
and AND2_1364 (wire937, n_476, n_426);
or OR2_1365 (wire938, n_475, n_431);
and AND2_1366 (wire941, wire940, n_476);
or OR2_1367 (n_487, wire942, n_475);
or OR2_1368 (n_492, wire943, n_474);
or OR2_1369 (n_496, wire944, n_473);
or OR2_1370 (wire947, wire946, n_471);
or OR2_1371 (n_498, wire948, n_470);
and AND2_1372 (wire952, n_466, n_465);
not NOT1_1373 (n_477, wire953);
or OR2_1374 (wire954, n_462, n_461);
not NOT1_1375 (n_480, wire955);
or OR2_1376 (wire956, n_458, n_457);
not NOT1_1377 (n_472, wire961);
and AND2_1378 (wire965, n_1564, n_423);
or OR2_1379 (wire982, n_1564, n_423);
not NOT1_1380 (n_434, wire987);
not NOT1_1381 (n_428, wire988);
and AND2_1382 (wire918, n_477, n_435);
or OR2_1383 (wire921, n_480, n_437);
or OR2_1384 (wire928, wire927, n_480);
and AND2_1385 (wire932, wire931, n_477);
not NOT1_1386 (n_486, wire933);
not NOT1_1387 (n_491, wire934);
not NOT1_1388 (n_495, wire935);
not NOT1_1389 (n_489, wire936);
not NOT1_1390 (n_493, wire937);
not NOT1_1391 (n_497, wire938);
or OR2_1392 (wire939, n_472, n_430);
not NOT1_1393 (n_508, wire941);
or OR2_1394 (n_488, wire945, n_472);
not NOT1_1395 (n_494, wire947);
not NOT1_1396 (n_484, wire952);
not NOT1_1397 (n_478, wire954);
not NOT1_1398 (n_481, wire956);
and AND2_1399 (wire969, wire968, n_428);
or OR2_1400 (n_456, wire974, n_434);
not NOT1_1401 (n_440, wire982);
not NOT1_1402 (wire1750, n_428);
and AND2_1403 (wire894, n_496, n_495);
and AND2_1404 (wire895, n_492, n_491);
and AND2_1405 (wire896, n_489, n_488);
and AND2_1406 (wire897, n_487, n_486);
or OR2_1407 (wire899, n_494, n_493);
and AND2_1408 (wire900, n_498, n_497);
or OR2_1409 (wire908, n_498, n_497);
or OR2_1410 (wire909, n_496, n_495);
and AND2_1411 (wire910, n_494, n_493);
or OR2_1412 (wire911, n_492, n_491);
or OR2_1413 (wire913, n_489, n_488);
or OR2_1414 (wire914, n_487, n_486);
or OR2_1415 (wire917, n_481, n_439);
not NOT1_1416 (n_506, wire918);
or OR2_1417 (wire919, n_478, n_436);
not NOT1_1418 (n_501, wire921);
and AND2_1419 (wire922, n_484, n_438);
and AND2_1420 (wire924, wire923, n_484);
or OR2_1421 (wire926, wire925, n_481);
not NOT1_1422 (n_505, wire928);
and AND2_1423 (wire929, n_456, n_455);
or OR2_1424 (n_502, wire930, n_478);
not NOT1_1425 (n_504, wire932);
not NOT1_1426 (n_500, wire939);
or OR2_1427 (wire957, n_456, n_455);
or OR2_1428 (wire966, wire965, n_440);
not NOT1_1429 (n_521, wire969);
or OR2_1430 (wire1751, wire1750, n_388);
and AND2_1431 (wire887, n_502, n_501);
or OR2_1432 (wire889, n_506, n_505);
and AND2_1433 (wire904, n_506, n_505);
or OR2_1434 (wire906, n_502, n_501);
not NOT1_1435 (n_513, wire908);
not NOT1_1436 (n_520, wire909);
not NOT1_1437 (n_514, wire910);
not NOT1_1438 (n_519, wire911);
not NOT1_1439 (n_518, wire913);
not NOT1_1440 (n_517, wire914);
not NOT1_1441 (n_503, wire917);
not NOT1_1442 (n_507, wire919);
not NOT1_1443 (n_510, wire922);
not NOT1_1444 (n2877, wire924);
not NOT1_1445 (n_509, wire926);
not NOT1_1446 (n_479, wire957);
not NOT1_1447 (n_468, wire966);
not NOT1_1448 (n_1563, wire1751);
or OR2_1449 (wire888, n_510, n_509);
and AND2_1450 (wire891, n_504, n_503);
and AND2_1451 (wire892, n_508, n_507);
or OR2_1452 (n_534, wire894, n_520);
or OR2_1453 (n_540, wire895, n_519);
or OR2_1454 (n_542, wire896, n_518);
or OR2_1455 (n_532, wire897, n_517);
and AND2_1456 (n_538, wire899, n_514);
or OR2_1457 (n_536, wire900, n_513);
and AND2_1458 (wire902, n_510, n_509);
or OR2_1459 (wire903, n_508, n_507);
not NOT1_1460 (n_526, wire904);
or OR2_1461 (wire905, n_504, n_503);
not NOT1_1462 (n_528, wire906);
and AND2_1463 (wire912, n_1563, n358);
or OR2_1464 (wire915, n_468, n_467);
or OR2_1465 (wire920, n_479, n_434);
or OR2_1466 (n_499, wire929, n_479);
or OR2_1467 (wire950, wire949, n_1563);
and AND2_1468 (wire951, n_468, n_467);
and AND2_1469 (wire853, n_536, n_535);
and AND2_1470 (wire861, n_540, n_539);
and AND2_1471 (wire862, n_542, n_541);
and AND2_1472 (wire863, n_534, n_533);
and AND2_1473 (wire865, n_532, n_531);
or OR2_1474 (wire868, n_538, n_537);
or OR2_1475 (wire878, n_542, n_541);
or OR2_1476 (wire879, n_540, n_539);
and AND2_1477 (wire880, n_538, n_537);
or OR2_1478 (wire881, n_536, n_535);
or OR2_1479 (wire883, n_534, n_533);
or OR2_1480 (wire884, n_532, n_531);
or OR2_1481 (n_545, wire887, n_528);
and AND2_1482 (n_553, wire889, n_526);
and AND2_1483 (wire890, n_500, n_499);
not NOT1_1484 (n_527, wire902);
not NOT1_1485 (n_523, wire903);
not NOT1_1486 (n_524, wire905);
or OR2_1487 (wire907, n_500, n_499);
not NOT1_1488 (n_512, wire920);
not NOT1_1489 (n_490, wire950);
not NOT1_1490 (n_482, wire951);
or OR2_1491 (wire844, n_553, n_552);
and AND2_1492 (wire846, n_545, n_544);
and AND2_1493 (wire871, n_553, n_552);
or OR2_1494 (wire875, n_545, n_544);
not NOT1_1495 (n_560, wire878);
not NOT1_1496 (n_561, wire879);
not NOT1_1497 (n_556, wire880);
not NOT1_1498 (n_564, wire881);
not NOT1_1499 (n_559, wire883);
not NOT1_1500 (n_558, wire884);
and AND2_1501 (n_551, wire888, n_527);
or OR2_1502 (n_547, wire891, n_524);
or OR2_1503 (n_555, wire892, n_523);
not NOT1_1504 (n_525, wire907);
or OR2_1505 (n_516, wire912, n_490);
and AND2_1506 (wire916, wire915, n_482);
not NOT1_1507 (wire1748, n_482);
or OR2_1508 (wire842, n_551, n_550);
and AND2_1509 (wire848, n_547, n_546);
and AND2_1510 (wire852, n_555, n_554);
or OR2_1511 (n_585, wire853, n_564);
or OR2_1512 (wire854, n_564, n_513);
or OR2_1513 (wire855, n_561, n_519);
or OR2_1514 (wire856, n_559, n_520);
or OR2_1515 (wire857, n_560, n_518);
or OR2_1516 (wire858, n_558, n_517);
and AND2_1517 (wire859, n_556, n_514);
or OR2_1518 (n_577, wire861, n_561);
or OR2_1519 (n_587, wire862, n_560);
or OR2_1520 (wire864, wire863, n_559);
or OR2_1521 (n_583, wire865, n_558);
and AND2_1522 (wire869, wire868, n_556);
or OR2_1523 (wire870, n_555, n_554);
not NOT1_1524 (n_571, wire871);
and AND2_1525 (wire872, n_551, n_550);
or OR2_1526 (wire874, n_547, n_546);
not NOT1_1527 (n_570, wire875);
and AND2_1528 (wire885, n_516, n_515);
or OR2_1529 (n_549, wire890, n_525);
or OR2_1530 (wire898, n_516, n_515);
not NOT1_1531 (n_511, wire916);
or OR2_1532 (wire1749, wire1748, n_440);
and AND2_1533 (wire837, n_571, n_526);
or OR2_1534 (wire841, n_570, n_528);
and AND2_1535 (wire845, wire844, n_571);
or OR2_1536 (wire847, wire846, n_570);
and AND2_1537 (wire851, n_549, n_548);
not NOT1_1538 (n_576, wire854);
not NOT1_1539 (n_586, wire855);
not NOT1_1540 (n_582, wire856);
not NOT1_1541 (n_597, wire857);
not NOT1_1542 (n_584, wire858);
not NOT1_1543 (n_580, wire859);
not NOT1_1544 (n_581, wire864);
not NOT1_1545 (n_591, wire869);
not NOT1_1546 (n_565, wire870);
not NOT1_1547 (n_572, wire872);
or OR2_1548 (wire873, n_549, n_548);
not NOT1_1549 (n_569, wire874);
and AND2_1550 (wire886, n_512, n_511);
not NOT1_1551 (n_530, wire898);
or OR2_1552 (wire901, n_512, n_511);
not NOT1_1553 (n_1562, wire1749);
or OR2_1554 (wire812, n_581, n_580);
and AND2_1555 (wire813, n_577, n_576);
and AND2_1556 (wire814, n_587, n_586);
and AND2_1557 (wire815, n_583, n_582);
and AND2_1558 (wire818, n_585, n_584);
or OR2_1559 (wire827, n_587, n_586);
or OR2_1560 (wire828, n_585, n_584);
or OR2_1561 (wire829, n_583, n_582);
and AND2_1562 (wire830, n_581, n_580);
or OR2_1563 (wire832, n_577, n_576);
or OR2_1564 (wire836, n_569, n_524);
not NOT1_1565 (n_588, wire837);
and AND2_1566 (wire838, n_572, n_527);
or OR2_1567 (wire839, n_565, n_523);
not NOT1_1568 (n_598, wire841);
and AND2_1569 (wire843, wire842, n_572);
not NOT1_1570 (n_593, wire845);
not NOT1_1571 (n_589, wire847);
or OR2_1572 (wire849, wire848, n_569);
or OR2_1573 (n_599, wire852, n_565);
not NOT1_1574 (n_566, wire873);
and AND2_1575 (wire876, n_1562, n_521);
or OR2_1576 (wire882, n_530, n_490);
or OR2_1577 (n_619, wire885, n_530);
or OR2_1578 (wire893, n_1562, n_521);
not NOT1_1579 (n_529, wire901);
and AND2_1580 (wire805, n_599, n_598);
or OR2_1581 (wire807, n_589, n_588);
or OR2_1582 (wire819, n_599, n_598);
and AND2_1583 (wire824, n_589, n_588);
not NOT1_1584 (n_606, wire827);
not NOT1_1585 (n_600, wire828);
not NOT1_1586 (n_605, wire829);
not NOT1_1587 (n_608, wire830);
not NOT1_1588 (n_607, wire832);
not NOT1_1589 (n_592, wire836);
not NOT1_1590 (n_594, wire838);
not NOT1_1591 (n_590, wire839);
or OR2_1592 (wire840, n_566, n_525);
not NOT1_1593 (n3211, wire843);
not NOT1_1594 (n_595, wire849);
or OR2_1595 (n_596, wire851, n_566);
not NOT1_1596 (n_557, wire882);
or OR2_1597 (n_563, wire886, n_529);
not NOT1_1598 (n_543, wire893);
or OR2_1599 (wire806, n_595, n_594);
and AND2_1600 (wire808, n_591, n_590);
and AND2_1601 (wire809, n_593, n_592);
and AND2_1602 (wire811, n_597, n_596);
and AND2_1603 (n_629, wire812, n_608);
or OR2_1604 (n_627, wire813, n_607);
or OR2_1605 (n_631, wire814, n_606);
or OR2_1606 (n_625, wire815, n_605);
or OR2_1607 (n_622, wire818, n_600);
not NOT1_1608 (n_618, wire819);
or OR2_1609 (wire820, n_597, n_596);
and AND2_1610 (wire821, n_595, n_594);
or OR2_1611 (wire822, n_593, n_592);
or OR2_1612 (wire823, n_591, n_590);
not NOT1_1613 (n_616, wire824);
and AND2_1614 (wire833, n_563, n_562);
and AND2_1615 (wire834, n_557, n375);
not NOT1_1616 (n_604, wire840);
or OR2_1617 (wire860, n_563, n_562);
or OR2_1618 (wire867, wire866, n_557);
or OR2_1619 (wire877, wire876, n_543);
or OR2_1620 (wire779, n_629, n_628);
and AND2_1621 (wire781, n_627, n_626);
and AND2_1622 (wire782, n_631, n_630);
and AND2_1623 (wire783, n_625, n_624);
and AND2_1624 (wire785, n_622, n_621);
or OR2_1625 (wire796, n_631, n_630);
and AND2_1626 (wire797, n_629, n_628);
or OR2_1627 (wire798, n_627, n_626);
or OR2_1628 (wire799, n_625, n_624);
or OR2_1629 (wire803, n_622, n_621);
or OR2_1630 (n_634, wire805, n_618);
and AND2_1631 (n_640, wire807, n_616);
not NOT1_1632 (n_609, wire820);
not NOT1_1633 (n_617, wire821);
not NOT1_1634 (n_612, wire822);
not NOT1_1635 (n_615, wire823);
not NOT1_1636 (n_575, wire860);
not NOT1_1637 (n_574, wire867);
not NOT1_1638 (n_568, wire877);
or OR2_1639 (wire755, n_640, n_639);
and AND2_1640 (wire771, n_634, n_633);
and AND2_1641 (wire791, n_640, n_639);
or OR2_1642 (wire794, n_634, n_633);
not NOT1_1643 (n_650, wire796);
not NOT1_1644 (n_652, wire797);
not NOT1_1645 (n_651, wire798);
not NOT1_1646 (n_649, wire799);
not NOT1_1647 (n_648, wire803);
and AND2_1648 (n_642, wire806, n_617);
or OR2_1649 (n_644, wire808, n_615);
or OR2_1650 (n_638, wire809, n_612);
or OR2_1651 (n_636, wire811, n_609);
or OR2_1652 (wire825, n_568, n_567);
or OR2_1653 (wire831, n_575, n_529);
or OR2_1654 (n_603, wire833, n_575);
or OR2_1655 (wire835, wire834, n_574);
and AND2_1656 (wire850, n_568, n_567);
or OR2_1657 (wire763, n_642, n_641);
and AND2_1658 (wire765, n_638, n_637);
and AND2_1659 (wire767, n_636, n_635);
and AND2_1660 (wire773, n_644, n_643);
and AND2_1661 (wire774, n_652, n_608);
or OR2_1662 (wire775, n_648, n_600);
or OR2_1663 (wire776, n_651, n_607);
or OR2_1664 (wire777, n_650, n_606);
or OR2_1665 (wire778, n_649, n_605);
and AND2_1666 (wire780, wire779, n_652);
or OR2_1667 (n_673, wire781, n_651);
or OR2_1668 (n_671, wire782, n_650);
or OR2_1669 (wire784, wire783, n_649);
or OR2_1670 (n_666, wire785, n_648);
or OR2_1671 (wire789, n_644, n_643);
and AND2_1672 (wire790, n_642, n_641);
not NOT1_1673 (n_662, wire791);
or OR2_1674 (wire792, n_638, n_637);
or OR2_1675 (wire793, n_636, n_635);
not NOT1_1676 (n_654, wire794);
and AND2_1677 (wire800, n_604, n_603);
or OR2_1678 (wire816, n_604, n_603);
not NOT1_1679 (n_611, wire831);
not NOT1_1680 (n_602, wire835);
not NOT1_1681 (n_578, wire850);
and AND2_1682 (wire756, wire755, n_662);
and AND2_1683 (wire757, n_662, n_616);
or OR2_1684 (wire762, n_654, n_618);
or OR2_1685 (wire772, wire771, n_654);
not NOT1_1686 (n_668, wire774);
not NOT1_1687 (n_672, wire775);
not NOT1_1688 (n_670, wire776);
not NOT1_1689 (n_685, wire777);
not NOT1_1690 (n_665, wire778);
not NOT1_1691 (n_683, wire780);
not NOT1_1692 (n_669, wire784);
not NOT1_1693 (n_653, wire789);
not NOT1_1694 (n_660, wire790);
not NOT1_1695 (n_659, wire792);
not NOT1_1696 (n_658, wire793);
or OR2_1697 (wire801, n_602, n_601);
not NOT1_1698 (n_623, wire816);
and AND2_1699 (wire817, n_602, n_601);
and AND2_1700 (wire826, wire825, n_578);
not NOT1_1701 (wire1746, n_578);
and AND2_1702 (wire732, n_673, n_672);
and AND2_1703 (wire733, n_671, n_670);
or OR2_1704 (wire734, n_669, n_668);
and AND2_1705 (wire735, n_666, n_665);
or OR2_1706 (wire748, n_673, n_672);
or OR2_1707 (wire749, n_671, n_670);
and AND2_1708 (wire750, n_669, n_668);
or OR2_1709 (wire753, n_666, n_665);
not NOT1_1710 (n_681, wire756);
not NOT1_1711 (n_686, wire757);
or OR2_1712 (wire758, n_653, n_615);
or OR2_1713 (wire759, n_658, n_609);
or OR2_1714 (wire760, n_659, n_612);
and AND2_1715 (wire761, n_660, n_617);
not NOT1_1716 (n_676, wire762);
and AND2_1717 (wire764, wire763, n_660);
or OR2_1718 (wire766, wire765, n_659);
or OR2_1719 (n_684, wire767, n_658);
not NOT1_1720 (n_687, wire772);
or OR2_1721 (n_677, wire773, n_653);
or OR2_1722 (n_647, wire800, n_623);
not NOT1_1723 (n_613, wire817);
not NOT1_1724 (n_610, wire826);
or OR2_1725 (wire1747, wire1746, n_543);
or OR2_1726 (wire726, n_687, n_686);
and AND2_1727 (wire727, n_685, n_684);
and AND2_1728 (wire730, n_677, n_676);
and AND2_1729 (wire740, n_687, n_686);
or OR2_1730 (wire741, n_685, n_684);
or OR2_1731 (wire745, n_677, n_676);
not NOT1_1732 (n_695, wire748);
not NOT1_1733 (n_694, wire749);
not NOT1_1734 (n_693, wire750);
and AND2_1735 (wire751, n_647, n_646);
not NOT1_1736 (n_692, wire753);
not NOT1_1737 (n_682, wire758);
not NOT1_1738 (n_690, wire759);
not NOT1_1739 (n_680, wire760);
not NOT1_1740 (n_688, wire761);
not NOT1_1741 (n3552, wire764);
not NOT1_1742 (n_689, wire766);
or OR2_1743 (wire786, n_647, n_646);
and AND2_1744 (wire795, n_611, n_610);
and AND2_1745 (wire802, wire801, n_613);
or OR2_1746 (wire810, n_611, n_610);
not NOT1_1747 (wire1744, n_613);
not NOT1_1748 (n_1561, wire1747);
and AND2_1749 (wire724, n_681, n_680);
and AND2_1750 (wire725, n_683, n_682);
or OR2_1751 (wire729, n_689, n_688);
or OR2_1752 (n_714, wire732, n_695);
or OR2_1753 (n_710, wire733, n_694);
and AND2_1754 (n_716, wire734, n_693);
or OR2_1755 (n_712, wire735, n_692);
and AND2_1756 (wire739, n_689, n_688);
not NOT1_1757 (n_703, wire740);
not NOT1_1758 (n_702, wire741);
or OR2_1759 (wire742, n_683, n_682);
or OR2_1760 (wire743, n_681, n_680);
not NOT1_1761 (n_698, wire745);
not NOT1_1762 (n_667, wire786);
and AND2_1763 (wire787, n_1561, n_619);
not NOT1_1764 (n_717, wire802);
or OR2_1765 (wire804, n_1561, n_619);
not NOT1_1766 (n_632, wire810);
or OR2_1767 (wire1745, wire1744, n_574);
or OR2_1768 (wire700, n_716, n_715);
and AND2_1769 (wire702, n_712, n_711);
and AND2_1770 (wire704, n_710, n_709);
and AND2_1771 (wire705, n_714, n_713);
and AND2_1772 (wire718, n_716, n_715);
or OR2_1773 (wire719, n_714, n_713);
or OR2_1774 (wire720, n_712, n_711);
or OR2_1775 (wire721, n_710, n_709);
and AND2_1776 (n_728, wire726, n_703);
or OR2_1777 (n_724, wire727, n_702);
or OR2_1778 (n_726, wire730, n_698);
not NOT1_1779 (n_699, wire739);
not NOT1_1780 (n_704, wire742);
not NOT1_1781 (n_705, wire743);
or OR2_1782 (n_691, wire751, n_667);
or OR2_1783 (wire752, n_667, n_623);
or OR2_1784 (n_657, wire795, n_632);
not NOT1_1785 (n_645, wire804);
not NOT1_1786 (n_1560, wire1745);
or OR2_1787 (wire684, n_728, n_727);
and AND2_1788 (wire688, n_724, n_723);
and AND2_1789 (wire689, n_726, n_725);
and AND2_1790 (wire710, n_728, n_727);
or OR2_1791 (wire711, n_726, n_725);
or OR2_1792 (wire712, n_724, n_723);
not NOT1_1793 (n_739, wire718);
not NOT1_1794 (n_736, wire719);
not NOT1_1795 (n_738, wire720);
not NOT1_1796 (n_737, wire721);
and AND2_1797 (wire722, n_691, n_690);
or OR2_1798 (n_721, wire724, n_705);
or OR2_1799 (n_732, wire725, n_704);
and AND2_1800 (n_730, wire729, n_699);
or OR2_1801 (wire736, n_691, n_690);
and AND2_1802 (wire746, n_1560, n392);
and AND2_1803 (wire747, n_657, n_656);
not NOT1_1804 (n_697, wire752);
or OR2_1805 (wire768, n_657, n_656);
or OR2_1806 (wire770, wire769, n_1560);
or OR2_1807 (wire788, wire787, n_645);
and AND2_1808 (wire675, n_732, n_731);
or OR2_1809 (wire682, n_730, n_729);
and AND2_1810 (wire686, n_721, n_720);
or OR2_1811 (wire696, n_736, n_695);
or OR2_1812 (wire697, n_738, n_692);
and AND2_1813 (wire698, n_739, n_693);
or OR2_1814 (wire699, n_737, n_694);
and AND2_1815 (wire701, wire700, n_739);
or OR2_1816 (wire703, wire702, n_738);
or OR2_1817 (n_759, wire704, n_737);
or OR2_1818 (n_755, wire705, n_736);
or OR2_1819 (wire708, n_732, n_731);
and AND2_1820 (wire709, n_730, n_729);
not NOT1_1821 (n_747, wire710);
not NOT1_1822 (n_744, wire711);
not NOT1_1823 (n_745, wire712);
or OR2_1824 (wire715, n_721, n_720);
not NOT1_1825 (n_708, wire736);
not NOT1_1826 (n_674, wire768);
not NOT1_1827 (n_675, wire770);
not NOT1_1828 (n_664, wire788);
and AND2_1829 (wire676, n_747, n_703);
or OR2_1830 (wire678, n_745, n_702);
or OR2_1831 (wire679, n_744, n_698);
and AND2_1832 (wire685, wire684, n_747);
or OR2_1833 (n_768, wire688, n_745);
or OR2_1834 (wire690, wire689, n_744);
not NOT1_1835 (n_758, wire696);
not NOT1_1836 (n_754, wire697);
not NOT1_1837 (n_757, wire698);
not NOT1_1838 (n_769, wire699);
not NOT1_1839 (n_775, wire701);
not NOT1_1840 (n_756, wire703);
not NOT1_1841 (n_750, wire708);
not NOT1_1842 (n_748, wire709);
not NOT1_1843 (n_746, wire715);
or OR2_1844 (n_735, wire722, n_708);
or OR2_1845 (wire737, n_664, n_663);
or OR2_1846 (wire744, n_674, n_632);
or OR2_1847 (n_701, wire746, n_675);
or OR2_1848 (n_696, wire747, n_674);
and AND2_1849 (wire754, n_664, n_663);
and AND2_1850 (wire647, n_769, n_768);
and AND2_1851 (wire652, n_755, n_754);
and AND2_1852 (wire653, n_759, n_758);
or OR2_1853 (wire654, n_757, n_756);
or OR2_1854 (wire661, n_769, n_768);
or OR2_1855 (wire669, n_759, n_758);
and AND2_1856 (wire670, n_757, n_756);
or OR2_1857 (wire671, n_755, n_754);
and AND2_1858 (wire673, n_735, n_734);
or OR2_1859 (n_767, wire675, n_750);
not NOT1_1860 (n_771, wire676);
or OR2_1861 (wire677, n_750, n_704);
not NOT1_1862 (n_778, wire678);
not NOT1_1863 (n_766, wire679);
and AND2_1864 (wire680, n_748, n_699);
or OR2_1865 (wire681, n_746, n_705);
and AND2_1866 (wire683, wire682, n_748);
not NOT1_1867 (n_764, wire685);
or OR2_1868 (wire687, wire686, n_746);
not NOT1_1869 (n_770, wire690);
or OR2_1870 (wire706, n_735, n_734);
and AND2_1871 (wire713, n_701, n_700);
and AND2_1872 (wire716, n_697, n_696);
or OR2_1873 (wire728, n_701, n_700);
or OR2_1874 (wire731, n_697, n_696);
not NOT1_1875 (n_707, wire744);
not NOT1_1876 (n_678, wire754);
and AND2_1877 (wire644, n_767, n_766);
or OR2_1878 (wire648, n_771, n_770);
and AND2_1879 (wire660, n_771, n_770);
not NOT1_1880 (n_787, wire661);
or OR2_1881 (wire662, n_767, n_766);
not NOT1_1882 (n_782, wire669);
not NOT1_1883 (n_781, wire670);
not NOT1_1884 (n_783, wire671);
not NOT1_1885 (n_774, wire677);
not NOT1_1886 (n_773, wire680);
not NOT1_1887 (n_763, wire681);
not NOT1_1888 (n3895, wire683);
not NOT1_1889 (n_772, wire687);
not NOT1_1890 (n_753, wire706);
not NOT1_1891 (n_722, wire728);
not NOT1_1892 (n_719, wire731);
and AND2_1893 (wire738, wire737, n_678);
not NOT1_1894 (wire1742, n_678);
and AND2_1895 (wire642, n_775, n_774);
or OR2_1896 (wire643, n_773, n_772);
and AND2_1897 (wire645, n_764, n_763);
or OR2_1898 (n_811, wire647, n_787);
or OR2_1899 (n_802, wire652, n_783);
or OR2_1900 (n_800, wire653, n_782);
and AND2_1901 (n_804, wire654, n_781);
or OR2_1902 (wire658, n_775, n_774);
and AND2_1903 (wire659, n_773, n_772);
not NOT1_1904 (n_786, wire660);
not NOT1_1905 (n_791, wire662);
or OR2_1906 (wire665, n_764, n_763);
or OR2_1907 (wire672, n_753, n_708);
or OR2_1908 (n_777, wire673, n_753);
or OR2_1909 (n_823, wire713, n_722);
or OR2_1910 (wire714, n_722, n_675);
or OR2_1911 (n_741, wire716, n_719);
not NOT1_1912 (n_706, wire738);
or OR2_1913 (wire1743, wire1742, n_645);
and AND2_1914 (wire602, n_811, n_810);
and AND2_1915 (wire616, n_800, n_799);
and AND2_1916 (wire617, n_802, n_801);
or OR2_1917 (wire619, n_804, n_803);
or OR2_1918 (wire633, n_811, n_810);
and AND2_1919 (wire637, n_804, n_803);
or OR2_1920 (wire638, n_802, n_801);
or OR2_1921 (wire639, n_800, n_799);
and AND2_1922 (wire641, n_778, n_777);
or OR2_1923 (n_813, wire644, n_791);
and AND2_1924 (n_817, wire648, n_786);
or OR2_1925 (wire656, n_778, n_777);
not NOT1_1926 (n_793, wire658);
not NOT1_1927 (n_792, wire659);
and AND2_1928 (wire663, n_741, n_740);
not NOT1_1929 (n_790, wire665);
not NOT1_1930 (n_785, wire672);
or OR2_1931 (wire695, n_741, n_740);
and AND2_1932 (wire707, n_707, n_706);
not NOT1_1933 (n_743, wire714);
or OR2_1934 (wire723, n_707, n_706);
not NOT1_1935 (n_1559, wire1743);
and AND2_1936 (wire600, n_813, n_812);
or OR2_1937 (wire606, n_817, n_816);
and AND2_1938 (wire628, n_817, n_816);
or OR2_1939 (wire630, n_813, n_812);
not NOT1_1940 (n_831, wire633);
not NOT1_1941 (n_820, wire637);
not NOT1_1942 (n_825, wire638);
not NOT1_1943 (n_821, wire639);
or OR2_1944 (n_819, wire642, n_793);
and AND2_1945 (n_815, wire643, n_792);
or OR2_1946 (n_809, wire645, n_790);
not NOT1_1947 (n_794, wire656);
and AND2_1948 (wire666, n_743, n409);
or OR2_1949 (wire692, wire691, n_743);
and AND2_1950 (wire693, n_1559, n_717);
not NOT1_1951 (n_765, wire695);
or OR2_1952 (wire717, n_1559, n_717);
not NOT1_1953 (n_733, wire723);
or OR2_1954 (wire598, n_815, n_814);
or OR2_1955 (n_859, wire602, n_831);
and AND2_1956 (wire608, n_809, n_808);
or OR2_1957 (wire612, n_831, n_787);
and AND2_1958 (wire614, n_819, n_818);
or OR2_1959 (n_840, wire616, n_821);
or OR2_1960 (wire618, wire617, n_825);
and AND2_1961 (wire620, wire619, n_820);
or OR2_1962 (wire622, n_825, n_783);
or OR2_1963 (wire625, n_821, n_782);
and AND2_1964 (wire626, n_820, n_781);
or OR2_1965 (wire627, n_819, n_818);
not NOT1_1966 (n_828, wire628);
and AND2_1967 (wire629, n_815, n_814);
not NOT1_1968 (n_833, wire630);
or OR2_1969 (wire634, n_809, n_808);
or OR2_1970 (n_827, wire641, n_794);
or OR2_1971 (n_784, wire663, n_765);
or OR2_1972 (wire664, n_765, n_719);
not NOT1_1973 (n_762, wire692);
or OR2_1974 (n_752, wire707, n_733);
not NOT1_1975 (n_742, wire717);
and AND2_1976 (wire597, n_827, n_826);
or OR2_1977 (wire601, wire600, n_833);
or OR2_1978 (wire605, n_833, n_791);
and AND2_1979 (wire607, wire606, n_828);
not NOT1_1980 (n_864, wire612);
and AND2_1981 (wire615, n_828, n_786);
not NOT1_1982 (n_842, wire618);
not NOT1_1983 (n_849, wire620);
or OR2_1984 (wire621, n_827, n_826);
not NOT1_1985 (n_839, wire622);
not NOT1_1986 (n_858, wire625);
not NOT1_1987 (n_841, wire626);
not NOT1_1988 (n_829, wire627);
not NOT1_1989 (n_832, wire629);
not NOT1_1990 (n_830, wire634);
and AND2_1991 (wire635, n_785, n_784);
or OR2_1992 (wire649, n_785, n_784);
and AND2_1993 (wire657, n_752, n_751);
not NOT1_1994 (n_796, wire664);
or OR2_1995 (wire667, wire666, n_762);
or OR2_1996 (wire674, n_752, n_751);
or OR2_1997 (wire694, wire693, n_742);
and AND2_1998 (wire569, n_859, n_858);
and AND2_1999 (wire574, n_840, n_839);
or OR2_2000 (wire575, n_842, n_841);
or OR2_2001 (wire581, n_859, n_858);
and AND2_2002 (wire595, n_842, n_841);
or OR2_2003 (wire596, n_840, n_839);
and AND2_2004 (wire599, wire598, n_832);
not NOT1_2005 (n_861, wire601);
not NOT1_2006 (n_850, wire605);
not NOT1_2007 (n_853, wire607);
or OR2_2008 (wire609, wire608, n_830);
and AND2_2009 (wire610, n_832, n_792);
or OR2_2010 (wire611, n_829, n_793);
or OR2_2011 (wire613, n_830, n_790);
or OR2_2012 (n_851, wire614, n_829);
not NOT1_2013 (n_860, wire615);
not NOT1_2014 (n_838, wire621);
not NOT1_2015 (n_807, wire649);
not NOT1_2016 (n_789, wire667);
not NOT1_2017 (n_776, wire674);
not NOT1_2018 (n_761, wire694);
or OR2_2019 (wire563, n_861, n_860);
and AND2_2020 (wire566, n_851, n_850);
and AND2_2021 (wire580, n_861, n_860);
not NOT1_2022 (n_871, wire581);
or OR2_2023 (wire585, n_851, n_850);
or OR2_2024 (wire594, n_838, n_794);
not NOT1_2025 (n_866, wire595);
not NOT1_2026 (n_867, wire596);
or OR2_2027 (n_863, wire597, n_838);
not NOT1_2028 (n4241, wire599);
not NOT1_2029 (n_855, wire609);
not NOT1_2030 (n_854, wire610);
not NOT1_2031 (n_848, wire611);
not NOT1_2032 (n_852, wire613);
or OR2_2033 (wire631, n_789, n_788);
or OR2_2034 (n_836, wire635, n_807);
and AND2_2035 (wire646, n_789, n_788);
or OR2_2036 (wire650, n_761, n_760);
or OR2_2037 (wire655, n_776, n_733);
or OR2_2038 (n_795, wire657, n_776);
and AND2_2039 (wire668, n_761, n_760);
and AND2_2040 (wire559, n_864, n_863);
and AND2_2041 (wire564, n_853, n_852);
or OR2_2042 (wire565, n_855, n_854);
and AND2_2043 (wire568, n_849, n_848);
or OR2_2044 (wire570, wire569, n_871);
or OR2_2045 (n_887, wire574, n_867);
and AND2_2046 (n_889, wire575, n_866);
or OR2_2047 (wire578, n_864, n_863);
not NOT1_2048 (n_878, wire580);
and AND2_2049 (wire583, n_855, n_854);
or OR2_2050 (wire584, n_853, n_852);
not NOT1_2051 (n_875, wire585);
or OR2_2052 (wire586, n_849, n_848);
and AND2_2053 (wire588, n_836, n_835);
not NOT1_2054 (n_873, wire594);
or OR2_2055 (wire603, n_836, n_835);
and AND2_2056 (wire624, n_796, n_795);
or OR2_2057 (wire640, n_796, n_795);
not NOT1_2058 (n_797, wire646);
not NOT1_2059 (n_806, wire655);
not NOT1_2060 (n_779, wire668);
and AND2_2061 (wire536, n_887, n_886);
or OR2_2062 (wire538, n_889, n_888);
and AND2_2063 (wire557, n_889, n_888);
or OR2_2064 (wire558, n_887, n_886);
and AND2_2065 (n_904, wire563, n_878);
or OR2_2066 (n_898, wire566, n_875);
not NOT1_2067 (n_896, wire570);
not NOT1_2068 (n_885, wire578);
not NOT1_2069 (n_876, wire583);
not NOT1_2070 (n_877, wire584);
not NOT1_2071 (n_872, wire586);
not NOT1_2072 (n_847, wire603);
and AND2_2073 (wire632, wire631, n_797);
not NOT1_2074 (n_822, wire640);
and AND2_2075 (wire651, wire650, n_779);
not NOT1_2076 (wire1738, n_797);
not NOT1_2077 (wire1740, n_779);
or OR2_2078 (wire521, n_904, n_903);
or OR2_2079 (wire525, n_896, n_895);
and AND2_2080 (wire532, n_898, n_897);
and AND2_2081 (wire546, n_904, n_903);
or OR2_2082 (wire549, n_898, n_897);
and AND2_2083 (wire550, n_896, n_895);
not NOT1_2084 (n_911, wire557);
not NOT1_2085 (n_912, wire558);
or OR2_2086 (wire560, wire559, n_885);
or OR2_2087 (n_894, wire564, n_877);
and AND2_2088 (n_900, wire565, n_876);
or OR2_2089 (n_902, wire568, n_872);
or OR2_2090 (wire587, n_847, n_807);
or OR2_2091 (n_874, wire588, n_847);
or OR2_2092 (n_846, wire624, n_822);
not NOT1_2093 (n_916, wire632);
not NOT1_2094 (n_805, wire651);
or OR2_2095 (wire1739, wire1738, n_762);
or OR2_2096 (wire1741, wire1740, n_742);
or OR2_2097 (wire514, n_900, n_899);
and AND2_2098 (wire523, n_894, n_893);
and AND2_2099 (wire527, n_902, n_901);
or OR2_2100 (wire534, n_912, n_867);
and AND2_2101 (wire535, n_911, n_866);
or OR2_2102 (wire537, wire536, n_912);
and AND2_2103 (wire539, wire538, n_911);
not NOT1_2104 (n_925, wire546);
or OR2_2105 (wire547, n_902, n_901);
and AND2_2106 (wire548, n_900, n_899);
not NOT1_2107 (n_915, wire549);
not NOT1_2108 (n_913, wire550);
or OR2_2109 (wire551, n_894, n_893);
and AND2_2110 (wire552, n_874, n_873);
not NOT1_2111 (n_909, wire560);
or OR2_2112 (wire567, n_874, n_873);
and AND2_2113 (wire576, n_846, n_845);
not NOT1_2114 (n_882, wire587);
or OR2_2115 (wire589, n_846, n_845);
and AND2_2116 (wire604, n_806, n_805);
or OR2_2117 (wire636, n_806, n_805);
not NOT1_2118 (n_1557, wire1739);
not NOT1_2119 (n_1558, wire1741);
or OR2_2120 (wire507, n_909, n_908);
or OR2_2121 (wire516, n_915, n_875);
and AND2_2122 (wire517, n_925, n_878);
and AND2_2123 (wire522, wire521, n_925);
and AND2_2124 (wire526, wire525, n_913);
or OR2_2125 (wire533, wire532, n_915);
not NOT1_2126 (n_943, wire534);
not NOT1_2127 (n_935, wire535);
not NOT1_2128 (n_934, wire537);
not NOT1_2129 (n_952, wire539);
and AND2_2130 (wire542, n_909, n_908);
not NOT1_2131 (n_921, wire547);
not NOT1_2132 (n_926, wire548);
not NOT1_2133 (n_922, wire551);
not NOT1_2134 (n_892, wire567);
and AND2_2135 (wire579, n_1557, n426);
not NOT1_2136 (n_865, wire589);
or OR2_2137 (wire591, wire590, n_1557);
and AND2_2138 (wire592, n_1558, n_823);
or OR2_2139 (wire623, n_1558, n_823);
not NOT1_2140 (n_834, wire636);
not NOT1_2141 (wire1734, n_913);
or OR2_2142 (wire487, n_935, n_934);
and AND2_2143 (wire506, n_935, n_934);
and AND2_2144 (wire515, wire514, n_926);
not NOT1_2145 (n_939, wire516);
not NOT1_2146 (n_948, wire517);
or OR2_2147 (wire518, n_921, n_872);
or OR2_2148 (wire519, n_922, n_877);
and AND2_2149 (wire520, n_926, n_876);
not NOT1_2150 (n_946, wire522);
or OR2_2151 (wire524, wire523, n_922);
not NOT1_2152 (n_944, wire526);
or OR2_2153 (n_940, wire527, n_921);
not NOT1_2154 (n_947, wire533);
not NOT1_2155 (n_923, wire542);
or OR2_2156 (wire553, wire552, n_892);
or OR2_2157 (n_881, wire576, n_865);
or OR2_2158 (wire577, n_865, n_822);
not NOT1_2159 (n_862, wire591);
or OR2_2160 (n_857, wire604, n_834);
not NOT1_2161 (n_843, wire623);
or OR2_2162 (wire1735, wire1734, n_871);
or OR2_2163 (wire477, n_948, n_947);
and AND2_2164 (wire480, n_940, n_939);
and AND2_2165 (wire485, n_944, n_943);
and AND2_2166 (wire497, n_948, n_947);
or OR2_2167 (wire499, n_944, n_943);
or OR2_2168 (wire502, n_940, n_939);
not NOT1_2169 (n_953, wire506);
and AND2_2170 (wire508, wire507, n_923);
not NOT1_2171 (n4591, wire515);
not NOT1_2172 (n_951, wire518);
not NOT1_2173 (n_945, wire519);
not NOT1_2174 (n_950, wire520);
not NOT1_2175 (n_949, wire524);
and AND2_2176 (wire543, n_882, n_881);
not NOT1_2177 (n_920, wire553);
or OR2_2178 (wire562, n_882, n_881);
and AND2_2179 (wire572, n_857, n_856);
not NOT1_2180 (n_891, wire577);
or OR2_2181 (n_884, wire579, n_862);
or OR2_2182 (wire582, n_857, n_856);
or OR2_2183 (wire593, wire592, n_843);
not NOT1_2184 (wire1732, n_923);
not NOT1_2185 (n_1555, wire1735);
and AND2_2186 (wire478, n_946, n_945);
and AND2_2187 (wire479, n_952, n_951);
or OR2_2188 (wire481, n_950, n_949);
and AND2_2189 (wire488, wire487, n_953);
or OR2_2190 (wire495, n_952, n_951);
and AND2_2191 (wire496, n_950, n_949);
not NOT1_2192 (n_973, wire497);
or OR2_2193 (wire498, n_946, n_945);
not NOT1_2194 (n_964, wire499);
or OR2_2195 (wire500, n_920, n_919);
not NOT1_2196 (n_970, wire502);
not NOT1_2197 (n_961, wire508);
and AND2_2198 (wire528, n_920, n_919);
and AND2_2199 (wire540, n_884, n_883);
or OR2_2200 (wire561, n_884, n_883);
not NOT1_2201 (n_907, wire562);
not NOT1_2202 (n_870, wire582);
not NOT1_2203 (n_869, wire593);
not NOT1_2204 (wire1726, n_953);
or OR2_2205 (wire1733, wire1732, n_885);
and AND2_2206 (wire472, n_961, n_1555);
and AND2_2207 (n_999, wire477, n_973);
or OR2_2208 (n_986, wire480, n_970);
or OR2_2209 (n_991, wire485, n_964);
not NOT1_2210 (n_982, wire488);
or OR2_2211 (wire489, n_961, n_1555);
not NOT1_2212 (n_971, wire495);
not NOT1_2213 (n_969, wire496);
not NOT1_2214 (n_972, wire498);
not NOT1_2215 (n_932, wire528);
or OR2_2216 (wire544, wire543, n_907);
or OR2_2217 (wire555, n_869, n_868);
not NOT1_2218 (n_910, wire561);
or OR2_2219 (wire571, n_870, n_834);
or OR2_2220 (n_890, wire572, n_870);
and AND2_2221 (wire573, n_869, n_868);
not NOT1_2222 (n_1554, wire1733);
and AND2_2223 (wire444, n_986, n_985);
or OR2_2224 (wire447, n_999, n_998);
and AND2_2225 (wire451, n_991, n_990);
and AND2_2226 (wire455, n_982, n_981);
and AND2_2227 (wire461, n_999, n_998);
or OR2_2228 (wire465, n_991, n_990);
or OR2_2229 (wire467, n_986, n_985);
or OR2_2230 (wire471, n_982, n_981);
or OR2_2231 (n_995, wire478, n_972);
or OR2_2232 (n_997, wire479, n_971);
and AND2_2233 (n_993, wire481, n_969);
not NOT1_2234 (n_980, wire489);
and AND2_2235 (wire501, wire500, n_932);
and AND2_2236 (wire529, n_891, n_890);
or OR2_2237 (n_1018, wire540, n_910);
or OR2_2238 (wire541, n_910, n_862);
not NOT1_2239 (n_931, wire544);
or OR2_2240 (wire554, n_891, n_890);
not NOT1_2241 (n_906, wire571);
not NOT1_2242 (n_879, wire573);
not NOT1_2243 (wire1730, n_932);
or OR2_2244 (wire436, n_993, n_992);
and AND2_2245 (wire449, n_995, n_994);
and AND2_2246 (wire452, n_997, n_996);
not NOT1_2247 (n_1012, wire461);
or OR2_2248 (wire462, n_997, n_996);
or OR2_2249 (wire463, n_995, n_994);
and AND2_2250 (wire464, n_993, n_992);
not NOT1_2251 (n_1010, wire465);
not NOT1_2252 (n_1015, wire467);
not NOT1_2253 (n_1005, wire471);
or OR2_2254 (n_1004, wire472, n_980);
or OR2_2255 (wire490, n_931, n_930);
not NOT1_2256 (n_965, wire501);
and AND2_2257 (wire509, n_931, n_930);
not NOT1_2258 (n_929, wire541);
not NOT1_2259 (n_918, wire554);
and AND2_2260 (wire556, wire555, n_879);
or OR2_2261 (wire1731, wire1730, n_892);
not NOT1_2262 (wire1736, n_879);
and AND2_2263 (wire432, n_1004, n_1003);
and AND2_2264 (wire438, n_1012, n_973);
or OR2_2265 (wire442, n_1010, n_964);
or OR2_2266 (wire443, n_1015, n_970);
or OR2_2267 (wire445, wire444, n_1015);
and AND2_2268 (wire448, wire447, n_1012);
or OR2_2269 (n_1036, wire451, n_1010);
or OR2_2270 (n_1040, wire455, n_1005);
or OR2_2271 (wire456, n_1004, n_1003);
not NOT1_2272 (n_1009, wire462);
not NOT1_2273 (n_1011, wire463);
not NOT1_2274 (n_1016, wire464);
and AND2_2275 (wire466, n_1554, n_965);
or OR2_2276 (wire482, n_1554, n_965);
and AND2_2277 (wire493, n_929, n443);
not NOT1_2278 (n_941, wire509);
or OR2_2279 (wire511, wire510, n_929);
or OR2_2280 (wire530, wire529, n_918);
not NOT1_2281 (n_905, wire556);
or OR2_2282 (wire1727, wire1726, n_1005);
not NOT1_2283 (n_1553, wire1731);
or OR2_2284 (wire1737, wire1736, n_843);
and AND2_2285 (wire437, wire436, n_1016);
not NOT1_2286 (n_1037, wire438);
and AND2_2287 (wire439, n_1016, n_969);
or OR2_2288 (wire440, n_1009, n_971);
or OR2_2289 (wire441, n_1011, n_972);
not NOT1_2290 (n_1045, wire442);
not NOT1_2291 (n_1031, wire443);
not NOT1_2292 (n_1038, wire445);
not NOT1_2293 (n_1030, wire448);
or OR2_2294 (wire450, wire449, n_1011);
or OR2_2295 (n_1032, wire452, n_1009);
not NOT1_2296 (n_1023, wire456);
not NOT1_2297 (n_987, wire482);
and AND2_2298 (wire491, wire490, n_941);
not NOT1_2299 (n_955, wire511);
and AND2_2300 (wire512, n_906, n_905);
not NOT1_2301 (n_938, wire530);
or OR2_2302 (wire545, n_906, n_905);
not NOT1_2303 (n_1551, wire1727);
not NOT1_2304 (wire1728, n_941);
not NOT1_2305 (n_1556, wire1737);
and AND2_2306 (wire402, n_1032, n_1031);
or OR2_2307 (wire405, n_1038, n_1037);
and AND2_2308 (wire406, n_1036, n_1551);
and AND2_2309 (wire420, n_1038, n_1037);
or OR2_2310 (wire421, n_1036, n_1551);
or OR2_2311 (wire423, n_1032, n_1031);
or OR2_2312 (wire431, n_1023, n_980);
or OR2_2313 (n_1046, wire432, n_1023);
not NOT1_2314 (n4946, wire437);
not NOT1_2315 (n_1034, wire439);
not NOT1_2316 (n_1039, wire440);
not NOT1_2317 (n_1029, wire441);
not NOT1_2318 (n_1033, wire450);
or OR2_2319 (n_1014, wire466, n_987);
or OR2_2320 (wire483, n_938, n_937);
not NOT1_2321 (n_975, wire491);
or OR2_2322 (wire494, wire493, n_955);
and AND2_2323 (wire503, n_938, n_937);
and AND2_2324 (wire504, n_1556, n_916);
or OR2_2325 (wire531, n_1556, n_916);
not NOT1_2326 (n_928, wire545);
or OR2_2327 (wire1729, wire1728, n_907);
and AND2_2328 (wire396, n_1046, n_1045);
and AND2_2329 (wire401, n_1040, n_1039);
or OR2_2330 (wire403, n_1034, n_1033);
and AND2_2331 (wire404, n_1030, n_1029);
or OR2_2332 (wire414, n_1046, n_1045);
or OR2_2333 (wire419, n_1040, n_1039);
not NOT1_2334 (n_1054, wire420);
not NOT1_2335 (n_1053, wire421);
and AND2_2336 (wire422, n_1034, n_1033);
not NOT1_2337 (n_1057, wire423);
or OR2_2338 (wire424, n_1030, n_1029);
and AND2_2339 (wire426, n_1014, n_1013);
not NOT1_2340 (n_1051, wire431);
or OR2_2341 (wire446, n_1014, n_1013);
and AND2_2342 (wire458, n_975, n_1553);
or OR2_2343 (wire474, n_975, n_1553);
not NOT1_2344 (n_979, wire494);
not NOT1_2345 (n_958, wire503);
or OR2_2346 (wire513, wire512, n_928);
not NOT1_2347 (n_936, wire531);
not NOT1_2348 (n_1552, wire1729);
or OR2_2349 (n_1076, wire402, n_1057);
and AND2_2350 (n_1084, wire405, n_1054);
or OR2_2351 (n_1078, wire406, n_1053);
not NOT1_2352 (n_1064, wire414);
not NOT1_2353 (n_1058, wire419);
not NOT1_2354 (n_1056, wire422);
not NOT1_2355 (n_1055, wire424);
not NOT1_2356 (n_1028, wire446);
or OR2_2357 (wire459, n_979, n_978);
and AND2_2358 (wire473, n_979, n_978);
not NOT1_2359 (n_1000, wire474);
and AND2_2360 (wire484, wire483, n_958);
or OR2_2361 (wire505, wire504, n_936);
not NOT1_2362 (n_957, wire513);
not NOT1_2363 (wire1724, n_958);
and AND2_2364 (wire370, n_1076, n_1075);
and AND2_2365 (wire372, n_1078, n_1077);
or OR2_2366 (wire378, n_1084, n_1083);
and AND2_2367 (wire385, n_1084, n_1083);
or OR2_2368 (wire388, n_1078, n_1077);
or OR2_2369 (wire389, n_1076, n_1075);
or OR2_2370 (n_1091, wire396, n_1064);
or OR2_2371 (n_1082, wire401, n_1058);
and AND2_2372 (n_1080, wire403, n_1056);
or OR2_2373 (n_1074, wire404, n_1055);
or OR2_2374 (wire425, n_1028, n_987);
or OR2_2375 (n_1052, wire426, n_1028);
or OR2_2376 (n_1022, wire458, n_1000);
not NOT1_2377 (n_988, wire473);
or OR2_2378 (wire475, n_957, n_956);
not NOT1_2379 (n_983, wire484);
and AND2_2380 (wire492, n_957, n_956);
not NOT1_2381 (n_963, wire505);
or OR2_2382 (wire1725, wire1724, n_918);
and AND2_2383 (wire355, n_1091, n_1090);
and AND2_2384 (wire365, n_1082, n_1081);
and AND2_2385 (wire366, n_1074, n_1073);
or OR2_2386 (wire368, n_1080, n_1079);
or OR2_2387 (wire380, n_1091, n_1090);
not NOT1_2388 (n_1092, wire385);
or OR2_2389 (wire386, n_1082, n_1081);
and AND2_2390 (wire387, n_1080, n_1079);
not NOT1_2391 (n_1098, wire388);
not NOT1_2392 (n_1099, wire389);
or OR2_2393 (wire390, n_1074, n_1073);
and AND2_2394 (wire395, n_1052, n_1051);
or OR2_2395 (wire407, n_1052, n_1051);
and AND2_2396 (wire415, n_1022, n_1021);
not NOT1_2397 (n_1063, wire425);
or OR2_2398 (wire433, n_1022, n_1021);
and AND2_2399 (wire453, n_1552, n_983);
and AND2_2400 (wire460, wire459, n_988);
or OR2_2401 (wire468, n_1552, n_983);
or OR2_2402 (wire469, n_963, n_962);
and AND2_2403 (wire486, n_963, n_962);
not NOT1_2404 (n_967, wire492);
not NOT1_2405 (wire1718, n_988);
not NOT1_2406 (n_1550, wire1725);
or OR2_2407 (wire359, n_1099, n_1057);
or OR2_2408 (wire362, n_1098, n_1053);
and AND2_2409 (wire364, n_1092, n_1054);
or OR2_2410 (wire371, wire370, n_1099);
or OR2_2411 (n_1125, wire372, n_1098);
and AND2_2412 (wire379, wire378, n_1092);
not NOT1_2413 (n_1109, wire380);
not NOT1_2414 (n_1103, wire386);
not NOT1_2415 (n_1100, wire387);
not NOT1_2416 (n_1102, wire390);
not NOT1_2417 (n_1065, wire407);
not NOT1_2418 (n_1044, wire433);
not NOT1_2419 (n_1110, wire460);
not NOT1_2420 (n_1008, wire468);
and AND2_2421 (wire476, wire475, n_967);
not NOT1_2422 (n_976, wire486);
or OR2_2423 (wire1719, wire1718, n_955);
not NOT1_2424 (wire1722, n_967);
or OR2_2425 (wire354, n_1109, n_1064);
or OR2_2426 (n_1132, wire355, n_1109);
not NOT1_2427 (n_1118, wire359);
and AND2_2428 (wire360, n_1100, n_1056);
or OR2_2429 (wire361, n_1103, n_1058);
not NOT1_2430 (n_1131, wire362);
or OR2_2431 (wire363, n_1102, n_1055);
not NOT1_2432 (n_1121, wire364);
or OR2_2433 (n_1119, wire365, n_1103);
or OR2_2434 (wire367, wire366, n_1102);
and AND2_2435 (wire369, wire368, n_1100);
not NOT1_2436 (n_1120, wire371);
not NOT1_2437 (n_1117, wire379);
or OR2_2438 (n_1097, wire395, n_1065);
or OR2_2439 (wire413, n_1044, n_1000);
or OR2_2440 (n_1062, wire415, n_1044);
or OR2_2441 (n_1027, wire453, n_1008);
and AND2_2442 (wire470, wire469, n_976);
not NOT1_2443 (n_1001, wire476);
not NOT1_2444 (n_1547, wire1719);
not NOT1_2445 (wire1720, n_976);
or OR2_2446 (wire1723, wire1722, n_928);
and AND2_2447 (wire317, n_1132, n_1131);
and AND2_2448 (wire331, n_1119, n_1118);
or OR2_2449 (wire332, n_1121, n_1120);
or OR2_2450 (wire337, n_1132, n_1131);
and AND2_2451 (wire346, n_1121, n_1120);
or OR2_2452 (wire347, n_1119, n_1118);
and AND2_2453 (wire350, n_1097, n_1096);
not NOT1_2454 (n_1141, wire354);
not NOT1_2455 (n_1123, wire360);
not NOT1_2456 (n_1124, wire361);
not NOT1_2457 (n_1116, wire363);
not NOT1_2458 (n_1122, wire367);
not NOT1_2459 (n5308, wire369);
or OR2_2460 (wire373, n_1097, n_1096);
and AND2_2461 (wire381, n_1063, n_1062);
or OR2_2462 (wire397, n_1063, n_1062);
and AND2_2463 (wire409, n_1027, n_1026);
and AND2_2464 (wire410, n_1547, n460);
not NOT1_2465 (n_1068, wire413);
or OR2_2466 (wire427, n_1027, n_1026);
or OR2_2467 (wire429, wire428, n_1547);
and AND2_2468 (wire434, n_1550, n_1001);
or OR2_2469 (wire457, n_1550, n_1001);
not NOT1_2470 (n_1006, wire470);
or OR2_2471 (wire1721, wire1720, n_936);
not NOT1_2472 (n_1549, wire1723);
and AND2_2473 (wire333, n_1117, n_1116);
or OR2_2474 (wire334, n_1123, n_1122);
and AND2_2475 (wire335, n_1125, n_1124);
not NOT1_2476 (n_1150, wire337);
or OR2_2477 (wire344, n_1125, n_1124);
and AND2_2478 (wire345, n_1123, n_1122);
not NOT1_2479 (n_1136, wire346);
not NOT1_2480 (n_1137, wire347);
or OR2_2481 (wire348, n_1117, n_1116);
not NOT1_2482 (n_1113, wire373);
not NOT1_2483 (n_1089, wire397);
not NOT1_2484 (n_1050, wire427);
not NOT1_2485 (n_1049, wire429);
and AND2_2486 (wire430, n_1549, n_1006);
or OR2_2487 (wire454, n_1549, n_1006);
not NOT1_2488 (n_1020, wire457);
not NOT1_2489 (n_1548, wire1721);
or OR2_2490 (wire318, wire317, n_1150);
or OR2_2491 (n_1156, wire331, n_1137);
and AND2_2492 (n_1154, wire332, n_1136);
not NOT1_2493 (n_1133, wire344);
not NOT1_2494 (n_1134, wire345);
not NOT1_2495 (n_1135, wire348);
or OR2_2496 (n_1142, wire350, n_1113);
or OR2_2497 (wire351, n_1113, n_1065);
or OR2_2498 (n_1108, wire381, n_1089);
or OR2_2499 (wire408, n_1050, n_1008);
or OR2_2500 (n_1067, wire409, n_1050);
or OR2_2501 (wire411, wire410, n_1049);
and AND2_2502 (wire417, n_1548, n_1018);
or OR2_2503 (n_1043, wire434, n_1020);
or OR2_2504 (wire435, n_1548, n_1018);
not NOT1_2505 (n_1024, wire454);
or OR2_2506 (wire289, n_1154, n_1153);
and AND2_2507 (wire296, n_1156, n_1155);
and AND2_2508 (wire308, n_1142, n_1141);
or OR2_2509 (wire314, n_1156, n_1155);
and AND2_2510 (wire315, n_1154, n_1153);
not NOT1_2511 (n_1169, wire318);
or OR2_2512 (wire327, n_1142, n_1141);
or OR2_2513 (n_1152, wire333, n_1135);
and AND2_2514 (n_1160, wire334, n_1134);
or OR2_2515 (wire336, wire335, n_1133);
and AND2_2516 (wire339, n_1108, n_1107);
not NOT1_2517 (n_1149, wire351);
or OR2_2518 (wire356, n_1108, n_1107);
and AND2_2519 (wire376, n_1068, n_1067);
or OR2_2520 (wire392, n_1068, n_1067);
and AND2_2521 (wire399, n_1043, n_1042);
not NOT1_2522 (n_1086, wire408);
not NOT1_2523 (n_1070, wire411);
or OR2_2524 (wire416, n_1043, n_1042);
or OR2_2525 (n_1048, wire430, n_1024);
not NOT1_2526 (n_1041, wire435);
or OR2_2527 (wire272, n_1169, n_1168);
or OR2_2528 (wire279, n_1160, n_1159);
and AND2_2529 (wire291, n_1152, n_1151);
and AND2_2530 (wire304, n_1169, n_1168);
and AND2_2531 (wire312, n_1160, n_1159);
not NOT1_2532 (n_1181, wire314);
not NOT1_2533 (n_1183, wire315);
or OR2_2534 (wire316, n_1152, n_1151);
not NOT1_2535 (n_1164, wire327);
not NOT1_2536 (n_1158, wire336);
not NOT1_2537 (n_1130, wire356);
or OR2_2538 (wire374, n_1070, n_1069);
and AND2_2539 (wire391, n_1070, n_1069);
not NOT1_2540 (n_1095, wire392);
and AND2_2541 (wire394, n_1048, n_1047);
or OR2_2542 (wire412, n_1048, n_1047);
not NOT1_2543 (n_1061, wire416);
or OR2_2544 (wire418, wire417, n_1041);
or OR2_2545 (wire285, n_1181, n_1137);
and AND2_2546 (wire288, n_1183, n_1136);
and AND2_2547 (wire290, wire289, n_1183);
or OR2_2548 (wire294, n_1158, n_1157);
or OR2_2549 (wire297, wire296, n_1181);
not NOT1_2550 (n_1184, wire304);
or OR2_2551 (wire309, wire308, n_1164);
not NOT1_2552 (n_1187, wire312);
and AND2_2553 (wire313, n_1158, n_1157);
not NOT1_2554 (n_1182, wire316);
or OR2_2555 (wire338, n_1130, n_1089);
or OR2_2556 (n_1148, wire339, n_1130);
or OR2_2557 (n_1115, wire376, n_1095);
not NOT1_2558 (n_1087, wire391);
or OR2_2559 (wire398, n_1061, n_1020);
or OR2_2560 (n_1085, wire399, n_1061);
not NOT1_2561 (n_1066, wire412);
not NOT1_2562 (n_1060, wire418);
and AND2_2563 (wire273, wire272, n_1184);
and AND2_2564 (wire280, wire279, n_1187);
and AND2_2565 (wire284, n_1187, n_1134);
not NOT1_2566 (n_1206, wire285);
not NOT1_2567 (n_1208, wire288);
not NOT1_2568 (n_1203, wire290);
or OR2_2569 (wire292, wire291, n_1182);
or OR2_2570 (wire293, n_1182, n_1135);
not NOT1_2571 (n_1209, wire297);
and AND2_2572 (wire301, n_1149, n_1148);
not NOT1_2573 (n_1180, wire309);
not NOT1_2574 (n_1172, wire313);
or OR2_2575 (wire319, n_1149, n_1148);
and AND2_2576 (wire325, n_1115, n_1114);
not NOT1_2577 (n_1166, wire338);
or OR2_2578 (wire349, n_1115, n_1114);
and AND2_2579 (wire357, n_1086, n_1085);
and AND2_2580 (wire375, wire374, n_1087);
or OR2_2581 (wire382, n_1060, n_1059);
or OR2_2582 (wire384, n_1086, n_1085);
or OR2_2583 (wire393, n_1066, n_1024);
or OR2_2584 (n_1093, wire394, n_1066);
not NOT1_2585 (n_1094, wire398);
and AND2_2586 (wire400, n_1060, n_1059);
not NOT1_2587 (wire1708, n_1184);
not NOT1_2588 (wire1714, n_1087);
or OR2_2589 (wire244, n_1209, n_1208);
and AND2_2590 (wire265, n_1209, n_1208);
or OR2_2591 (wire267, n_1180, n_1179);
not NOT1_2592 (n_1222, wire273);
not NOT1_2593 (n5672, wire280);
not NOT1_2594 (n_1213, wire284);
not NOT1_2595 (n_1214, wire292);
not NOT1_2596 (n_1202, wire293);
and AND2_2597 (wire295, wire294, n_1172);
and AND2_2598 (wire298, n_1180, n_1179);
not NOT1_2599 (n_1174, wire319);
not NOT1_2600 (n_1143, wire349);
and AND2_2601 (wire352, n_1094, n_1093);
not NOT1_2602 (n_1219, wire375);
or OR2_2603 (wire377, n_1094, n_1093);
not NOT1_2604 (n_1106, wire384);
not NOT1_2605 (n_1105, wire393);
not NOT1_2606 (n_1071, wire400);
or OR2_2607 (wire1709, wire1708, n_1150);
not NOT1_2608 (wire1710, n_1172);
or OR2_2609 (wire1715, wire1714, n_1049);
and AND2_2610 (wire240, n_1203, n_1202);
or OR2_2611 (wire241, n_1214, n_1213);
and AND2_2612 (wire261, n_1214, n_1213);
not NOT1_2613 (n_1224, wire265);
or OR2_2614 (wire269, n_1203, n_1202);
not NOT1_2615 (n_1207, wire295);
not NOT1_2616 (n_1196, wire298);
or OR2_2617 (wire302, wire301, n_1174);
or OR2_2618 (n_1165, wire325, n_1143);
or OR2_2619 (wire326, n_1143, n_1095);
or OR2_2620 (n_1129, wire357, n_1106);
not NOT1_2621 (n_1112, wire377);
and AND2_2622 (wire383, wire382, n_1071);
not NOT1_2623 (n_1542, wire1709);
or OR2_2624 (wire1711, wire1710, n_1133);
not NOT1_2625 (n_1545, wire1715);
not NOT1_2626 (wire1716, n_1071);
and AND2_2627 (wire245, wire244, n_1224);
and AND2_2628 (wire246, n_1207, n_1206);
not NOT1_2629 (n_1235, wire261);
or OR2_2630 (wire266, n_1207, n_1206);
and AND2_2631 (wire268, wire267, n_1196);
not NOT1_2632 (n_1236, wire269);
and AND2_2633 (wire286, n_1166, n_1165);
not NOT1_2634 (n_1195, wire302);
or OR2_2635 (wire307, n_1166, n_1165);
and AND2_2636 (wire321, n_1129, n_1128);
and AND2_2637 (wire322, n_1545, n477);
not NOT1_2638 (n_1178, wire326);
or OR2_2639 (wire340, n_1129, n_1128);
or OR2_2640 (wire342, wire341, n_1545);
or OR2_2641 (n_1140, wire352, n_1112);
not NOT1_2642 (n_1104, wire383);
not NOT1_2643 (wire1698, n_1224);
not NOT1_2644 (wire1704, n_1196);
not NOT1_2645 (n_1543, wire1711);
or OR2_2646 (wire1717, wire1716, n_1041);
and AND2_2647 (wire235, n_1222, n_1543);
or OR2_2648 (n_1254, wire240, n_1236);
and AND2_2649 (n_1260, wire241, n_1235);
not NOT1_2650 (n_1256, wire245);
or OR2_2651 (wire256, n_1222, n_1543);
or OR2_2652 (wire259, n_1195, n_1194);
not NOT1_2653 (n_1233, wire266);
not NOT1_2654 (n_1230, wire268);
and AND2_2655 (wire274, n_1195, n_1194);
not NOT1_2656 (n_1186, wire307);
and AND2_2657 (wire310, n_1140, n_1139);
or OR2_2658 (wire328, n_1140, n_1139);
not NOT1_2659 (n_1147, wire340);
not NOT1_2660 (n_1146, wire342);
and AND2_2661 (wire343, n_1105, n_1104);
or OR2_2662 (wire358, n_1105, n_1104);
or OR2_2663 (wire1705, wire1704, n_1164);
not NOT1_2664 (n_1546, wire1717);
and AND2_2665 (wire203, n_1256, n_1255);
and AND2_2666 (wire204, n_1254, n_1253);
or OR2_2667 (wire209, n_1260, n_1259);
and AND2_2668 (wire222, n_1260, n_1259);
or OR2_2669 (wire224, n_1256, n_1255);
or OR2_2670 (wire225, n_1254, n_1253);
and AND2_2671 (wire226, n_1230, n_1542);
or OR2_2672 (wire247, wire246, n_1233);
or OR2_2673 (wire250, n_1230, n_1542);
not NOT1_2674 (n_1243, wire256);
not NOT1_2675 (n_1204, wire274);
or OR2_2676 (wire287, wire286, n_1186);
or OR2_2677 (wire320, n_1147, n_1106);
or OR2_2678 (n_1177, wire321, n_1147);
or OR2_2679 (wire323, wire322, n_1146);
not NOT1_2680 (n_1163, wire328);
and AND2_2681 (wire329, n_1546, n_1110);
or OR2_2682 (wire353, n_1546, n_1110);
not NOT1_2683 (n_1126, wire358);
not NOT1_2684 (n_1540, wire1705);
not NOT1_2685 (n_1277, wire222);
not NOT1_2686 (n_1282, wire224);
not NOT1_2687 (n_1281, wire225);
or OR2_2688 (n_1269, wire235, n_1243);
not NOT1_2689 (n_1258, wire247);
not NOT1_2690 (n_1252, wire250);
and AND2_2691 (wire260, wire259, n_1204);
and AND2_2692 (wire277, n_1177, n_1178);
not NOT1_2693 (n_1201, wire287);
or OR2_2694 (wire299, n_1178, n_1177);
or OR2_2695 (wire306, n_1163, n_1112);
or OR2_2696 (n_1188, wire310, n_1163);
not NOT1_2697 (n_1189, wire320);
not NOT1_2698 (n_1176, wire323);
or OR2_2699 (n_1145, wire343, n_1126);
not NOT1_2700 (n_1138, wire353);
not NOT1_2701 (wire1702, n_1204);
and AND2_2702 (wire194, n_1269, n_1268);
and AND2_2703 (wire202, n_1277, n_1235);
or OR2_2704 (n_1303, wire203, n_1282);
or OR2_2705 (wire205, wire204, n_1281);
or OR2_2706 (wire206, n_1258, n_1257);
or OR2_2707 (wire208, n_1281, n_1236);
and AND2_2708 (wire210, wire209, n_1277);
or OR2_2709 (wire216, n_1269, n_1268);
and AND2_2710 (wire223, n_1258, n_1257);
or OR2_2711 (n_1284, wire226, n_1252);
or OR2_2712 (wire248, n_1201, n_1200);
not NOT1_2713 (n_1242, wire260);
and AND2_2714 (wire263, n_1189, n_1188);
and AND2_2715 (wire270, n_1201, n_1200);
or OR2_2716 (wire275, n_1176, n_1175);
or OR2_2717 (wire281, n_1189, n_1188);
not NOT1_2718 (n_1193, wire299);
and AND2_2719 (wire300, n_1176, n_1175);
and AND2_2720 (wire305, n_1145, n_1144);
not NOT1_2721 (n_1199, wire306);
or OR2_2722 (wire324, n_1145, n_1144);
or OR2_2723 (wire330, wire329, n_1138);
or OR2_2724 (wire1699, wire1698, n_1282);
or OR2_2725 (wire1703, wire1702, n_1174);
and AND2_2726 (wire184, n_1284, n_1283);
or OR2_2727 (wire201, n_1284, n_1283);
not NOT1_2728 (n_1298, wire202);
not NOT1_2729 (n_1299, wire205);
not NOT1_2730 (n_1302, wire208);
not NOT1_2731 (n5971, wire210);
not NOT1_2732 (n_1292, wire216);
and AND2_2733 (wire217, n_1242, n_1540);
not NOT1_2734 (n_1270, wire223);
or OR2_2735 (wire236, n_1242, n_1540);
not NOT1_2736 (n_1217, wire270);
or OR2_2737 (wire278, wire277, n_1193);
not NOT1_2738 (n_1210, wire281);
not NOT1_2739 (n_1191, wire300);
not NOT1_2740 (n_1167, wire324);
not NOT1_2741 (n_1162, wire330);
not NOT1_2742 (n_1537, wire1699);
not NOT1_2743 (n_1539, wire1703);
or OR2_2744 (wire173, n_1299, n_1298);
and AND2_2745 (wire175, n_1303, n_1302);
or OR2_2746 (wire186, n_1303, n_1302);
and AND2_2747 (wire190, n_1299, n_1298);
or OR2_2748 (n_1306, wire194, n_1292);
or OR2_2749 (wire195, n_1292, n_1243);
not NOT1_2750 (n_1304, wire201);
and AND2_2751 (wire207, wire206, n_1270);
not NOT1_2752 (n_1267, wire236);
and AND2_2753 (wire249, wire248, n_1217);
or OR2_2754 (wire264, wire263, n_1210);
and AND2_2755 (wire276, wire275, n_1191);
not NOT1_2756 (n_1216, wire278);
or OR2_2757 (wire282, n_1162, n_1161);
or OR2_2758 (wire303, n_1167, n_1126);
or OR2_2759 (n_1198, wire305, n_1167);
and AND2_2760 (wire311, n_1162, n_1161);
not NOT1_2761 (wire1688, n_1270);
not NOT1_2762 (wire1700, n_1217);
not NOT1_2763 (wire1706, n_1191);
or OR2_2764 (n_1314, wire184, n_1304);
or OR2_2765 (wire185, n_1304, n_1252);
not NOT1_2766 (n_1316, wire186);
not NOT1_2767 (n_1317, wire190);
not NOT1_2768 (n_1313, wire195);
not NOT1_2769 (n_1294, wire207);
or OR2_2770 (n_1291, wire217, n_1267);
or OR2_2771 (wire238, n_1216, n_1215);
not NOT1_2772 (n_1247, wire249);
and AND2_2773 (wire254, n_1199, n_1198);
and AND2_2774 (wire258, n_1216, n_1215);
not NOT1_2775 (n_1228, wire264);
or OR2_2776 (wire271, n_1199, n_1198);
not NOT1_2777 (n_1318, wire276);
not NOT1_2778 (n_1212, wire303);
not NOT1_2779 (n_1170, wire311);
or OR2_2780 (wire1689, wire1688, n_1233);
or OR2_2781 (wire1701, wire1700, n_1186);
or OR2_2782 (wire1707, wire1706, n_1146);
and AND2_2783 (wire159, n_1314, n_1313);
and AND2_2784 (wire174, wire173, n_1317);
or OR2_2785 (n_1337, wire175, n_1316);
and AND2_2786 (wire176, n_1294, n_1537);
or OR2_2787 (wire177, n_1314, n_1313);
and AND2_2788 (wire179, n_1291, n_1290);
not NOT1_2789 (n_1324, wire185);
or OR2_2790 (wire193, n_1294, n_1537);
or OR2_2791 (wire196, n_1291, n_1290);
and AND2_2792 (wire215, n_1539, n_1247);
or OR2_2793 (wire227, n_1228, n_1227);
or OR2_2794 (wire231, n_1539, n_1247);
and AND2_2795 (wire251, n_1228, n_1227);
not NOT1_2796 (n_1231, wire258);
not NOT1_2797 (n_1223, wire271);
and AND2_2798 (wire283, wire282, n_1170);
not NOT1_2799 (n_1532, wire1689);
not NOT1_2800 (n_1538, wire1701);
not NOT1_2801 (n_1541, wire1707);
not NOT1_2802 (wire1712, n_1170);
and AND2_2803 (wire134, n_1337, n_1336);
or OR2_2804 (wire156, n_1337, n_1336);
and AND2_2805 (wire165, n_1306, n_1532);
not NOT1_2806 (n_1328, wire174);
not NOT1_2807 (n_1334, wire177);
or OR2_2808 (wire183, n_1306, n_1532);
not NOT1_2809 (n_1315, wire193);
not NOT1_2810 (n_1312, wire196);
and AND2_2811 (wire229, n_1541, n494);
not NOT1_2812 (n_1272, wire231);
and AND2_2813 (wire239, wire238, n_1231);
not NOT1_2814 (n_1239, wire251);
or OR2_2815 (wire253, wire252, n_1541);
or OR2_2816 (wire255, wire254, n_1223);
not NOT1_2817 (n_1211, wire283);
not NOT1_2818 (wire1696, n_1231);
or OR2_2819 (wire1713, wire1712, n_1138);
not NOT1_2820 (n_1363, wire156);
or OR2_2821 (n_1359, wire159, n_1334);
or OR2_2822 (n_1339, wire176, n_1315);
or OR2_2823 (wire178, n_1312, n_1267);
or OR2_2824 (n_1325, wire179, n_1312);
not NOT1_2825 (n_1327, wire183);
or OR2_2826 (n_1301, wire215, n_1272);
and AND2_2827 (wire228, wire227, n_1239);
not NOT1_2828 (n_1266, wire239);
and AND2_2829 (wire242, n_1212, n_1211);
not NOT1_2830 (n_1249, wire253);
not NOT1_2831 (n_1238, wire255);
or OR2_2832 (wire262, n_1212, n_1211);
not NOT1_2833 (wire1682, n_1328);
not NOT1_2834 (wire1694, n_1239);
or OR2_2835 (wire1697, wire1696, n_1193);
not NOT1_2836 (n_1544, wire1713);
and AND2_2837 (wire1759, wire1758, n_1328);
and AND2_2838 (wire116, n_1359, n_1358);
and AND2_2839 (wire133, n_1339, n_1338);
or OR2_2840 (wire135, wire134, n_1363);
or OR2_2841 (wire137, n_1363, n_1316);
or OR2_2842 (wire140, n_1359, n_1358);
and AND2_2843 (wire148, n_1325, n_1324);
or OR2_2844 (wire155, n_1339, n_1338);
or OR2_2845 (n_1349, wire165, n_1327);
or OR2_2846 (wire167, n_1325, n_1324);
and AND2_2847 (wire169, n_1301, n_1300);
not NOT1_2848 (n_1344, wire178);
or OR2_2849 (wire187, n_1301, n_1300);
and AND2_2850 (wire198, n_1266, n_1538);
or OR2_2851 (wire218, n_1266, n_1538);
or OR2_2852 (wire220, n_1238, n_1237);
not NOT1_2853 (n_1275, wire228);
or OR2_2854 (wire230, wire229, n_1249);
and AND2_2855 (wire233, n_1544, n_1219);
and AND2_2856 (wire237, n_1238, n_1237);
or OR2_2857 (wire257, n_1544, n_1219);
not NOT1_2858 (n_1234, wire262);
and AND2_2859 (wire1683, wire1682, n_34);
or OR2_2860 (wire1695, wire1694, n_1210);
not NOT1_2861 (n_1536, wire1697);
not NOT1_2862 (n_1567, wire1759);
and AND2_2863 (wire126, n_1349, n_1348);
not NOT1_2864 (n_1388, wire135);
not NOT1_2865 (n_1378, wire137);
not NOT1_2866 (n_1380, wire140);
or OR2_2867 (wire149, n_1349, n_1348);
not NOT1_2868 (n_1357, wire155);
not NOT1_2869 (n_1350, wire167);
not NOT1_2870 (n_1321, wire187);
and AND2_2871 (wire192, n_1536, n_1275);
or OR2_2872 (wire213, n_1536, n_1275);
not NOT1_2873 (n_1285, wire218);
not NOT1_2874 (n_1274, wire230);
not NOT1_2875 (n_1250, wire237);
or OR2_2876 (wire243, wire242, n_1234);
not NOT1_2877 (n_1244, wire257);
not NOT1_2878 (n_1529, wire1683);
not NOT1_2879 (n_1535, wire1695);
or OR2_2880 (n_1399, wire116, n_1380);
and AND2_2881 (wire117, n_1529, n_1567);
or OR2_2882 (wire120, n_1380, n_1334);
and AND2_2883 (wire127, n_1529, n_1317);
or OR2_2884 (n_1379, wire133, n_1357);
or OR2_2885 (wire141, n_1357, n_1315);
or OR2_2886 (n_1370, wire148, n_1350);
not NOT1_2887 (n_1373, wire149);
or OR2_2888 (n_1343, wire169, n_1321);
or OR2_2889 (wire170, n_1321, n_1272);
or OR2_2890 (wire188, n_1274, n_1273);
or OR2_2891 (n_1311, wire198, n_1285);
not NOT1_2892 (n_1295, wire213);
and AND2_2893 (wire214, n_1274, n_1273);
and AND2_2894 (wire221, wire220, n_1250);
or OR2_2895 (wire234, wire233, n_1244);
not NOT1_2896 (n_1246, wire243);
not NOT1_2897 (wire1692, n_1250);
and AND2_2898 (wire99, n_1379, n_1378);
and AND2_2899 (wire104, n_1370, n_1369);
or OR2_2900 (wire118, wire117, n_373);
not NOT1_2901 (n_1408, wire120);
or OR2_2902 (wire121, n_1379, n_1378);
or OR2_2903 (wire124, n_1373, n_1327);
or OR2_2904 (n_1394, wire126, n_1373);
not NOT1_2905 (n_1387, wire127);
or OR2_2906 (wire129, n_1370, n_1369);
and AND2_2907 (wire138, n_1344, n_1343);
not NOT1_2908 (n_1393, wire141);
or OR2_2909 (wire153, n_1344, n_1343);
and AND2_2910 (wire161, n_1311, n_1310);
not NOT1_2911 (n_1347, wire170);
or OR2_2912 (wire180, n_1311, n_1310);
or OR2_2913 (n_1323, wire192, n_1295);
or OR2_2914 (wire211, n_1246, n_1245);
not NOT1_2915 (n_1288, wire214);
not NOT1_2916 (n_1286, wire221);
and AND2_2917 (wire232, n_1246, n_1245);
not NOT1_2918 (n_1262, wire234);
or OR2_2919 (wire1693, wire1692, n_1223);
and AND2_2920 (wire84, n_1387, n_1388);
and AND2_2921 (wire94, n_1394, n_1393);
or OR2_2922 (wire106, n_1394, n_1393);
or OR2_2923 (wire112, n_1388, n_1387);
not NOT1_2924 (n_1413, wire118);
not NOT1_2925 (n_1403, wire121);
not NOT1_2926 (n_1398, wire124);
not NOT1_2927 (n_1392, wire129);
and AND2_2928 (wire151, n_1323, n_1322);
not NOT1_2929 (n_1362, wire153);
or OR2_2930 (wire168, n_1323, n_1322);
not NOT1_2931 (n_1331, wire180);
and AND2_2932 (wire182, n_1535, n_1286);
and AND2_2933 (wire189, wire188, n_1288);
or OR2_2934 (wire197, n_1535, n_1286);
or OR2_2935 (wire199, n_1262, n_1261);
and AND2_2936 (wire219, n_1262, n_1261);
not NOT1_2937 (n_1263, wire232);
not NOT1_2938 (wire1684, n_1288);
not NOT1_2939 (n_1534, wire1693);
and AND2_2940 (wire83, n_1399, n_1398);
or OR2_2941 (wire89, n_1413, n_1412);
and AND2_2942 (wire90, n_1413, n_1412);
or OR2_2943 (n_1422, wire99, n_1403);
or OR2_2944 (wire102, n_1399, n_1398);
or OR2_2945 (n_1409, wire104, n_1392);
not NOT1_2946 (n_1410, wire106);
or OR2_2947 (wire109, n_1392, n_1350);
not NOT1_2948 (n_1421, wire112);
or OR2_2949 (n_1386, wire138, n_1362);
or OR2_2950 (n_1346, wire161, n_1331);
or OR2_2951 (wire162, n_1331, n_1285);
not NOT1_2952 (n_1345, wire168);
not NOT1_2953 (n_1417, wire189);
not NOT1_2954 (n_1307, wire197);
and AND2_2955 (wire212, wire211, n_1263);
not NOT1_2956 (n_1279, wire219);
or OR2_2957 (wire1685, wire1684, n_1249);
not NOT1_2958 (wire1690, n_1263);
and AND2_2959 (wire64, n_1422, n_1421);
and AND2_2960 (wire74, n_1409, n_1408);
or OR2_2961 (wire80, n_1422, n_1421);
or OR2_2962 (wire85, wire84, n_1421);
not NOT1_2963 (wire91, wire90);
or OR2_2964 (n_1456, wire94, n_1410);
or OR2_2965 (wire95, n_1409, n_1408);
and AND2_2966 (wire98, n_1386, n_1385);
not NOT1_2967 (n_1419, wire102);
not NOT1_2968 (n_1428, wire109);
or OR2_2969 (wire113, n_1386, n_1385);
and AND2_2970 (wire128, n_1347, n_1346);
or OR2_2971 (wire150, n_1347, n_1346);
or OR2_2972 (n_1355, wire151, n_1345);
or OR2_2973 (wire152, n_1345, n_1295);
not NOT1_2974 (n_1356, wire162);
or OR2_2975 (n_1333, wire182, n_1307);
and AND2_2976 (wire200, wire199, n_1279);
not NOT1_2977 (n_1296, wire212);
not NOT1_2978 (n_1530, wire1685);
not NOT1_2979 (wire1686, n_1279);
or OR2_2980 (wire1691, wire1690, n_1234);
not NOT1_2981 (n_1436, wire80);
or OR2_2982 (n_1470, wire83, n_1419);
not NOT1_2983 (n6150, wire85);
and AND2_2984 (wire92, wire91, wire89);
not NOT1_2985 (n_1429, wire95);
not NOT1_2986 (n_1397, wire113);
and AND2_2987 (wire122, n_1356, n_1355);
or OR2_2988 (wire142, n_1356, n_1355);
and AND2_2989 (wire143, n_1530, n511);
and AND2_2990 (wire145, n_1333, n_1332);
not NOT1_2991 (n_1371, wire150);
not NOT1_2992 (n_1366, wire152);
or OR2_2993 (wire160, n_1333, n_1332);
or OR2_2994 (wire164, wire163, n_1530);
and AND2_2995 (wire171, n_1534, n_1296);
or OR2_2996 (wire191, n_1534, n_1296);
not NOT1_2997 (n_1308, wire200);
or OR2_2998 (wire1687, wire1686, n_1244);
not NOT1_2999 (n_1533, wire1691);
or OR2_3000 (n6160, wire64, n_1436);
or OR2_3001 (wire67, n_1436, n_1403);
or OR2_3002 (n_1479, wire74, n_1429);
not NOT1_3003 (n6123, wire92);
or OR2_3004 (n_1427, wire98, n_1397);
or OR2_3005 (wire103, n_1397, n_1362);
or OR2_3006 (n_1391, wire128, n_1371);
not NOT1_3007 (n_1377, wire142);
not NOT1_3008 (n_1353, wire160);
not NOT1_3009 (n_1354, wire164);
and AND2_3010 (wire166, n_1533, n_1308);
or OR2_3011 (wire181, n_1533, n_1308);
not NOT1_3012 (n_1320, wire191);
not NOT1_3013 (n_1531, wire1687);
and AND2_3014 (wire62, n_1428, n_1427);
not NOT1_3015 (n_1457, wire67);
or OR2_3016 (wire75, n_1428, n_1427);
and AND2_3017 (wire88, n_1391, n_1390);
not NOT1_3018 (n_1431, wire103);
or OR2_3019 (wire110, n_1391, n_1390);
or OR2_3020 (n_1405, wire122, n_1377);
or OR2_3021 (wire144, wire143, n_1354);
or OR2_3022 (n_1365, wire145, n_1353);
or OR2_3023 (wire146, n_1353, n_1307);
and AND2_3024 (wire157, n_1531, n_1318);
or OR2_3025 (n_1342, wire171, n_1320);
or OR2_3026 (wire172, n_1531, n_1318);
not NOT1_3027 (n_1326, wire181);
and AND2_3028 (wire42, n_1457, n_1456);
or OR2_3029 (wire52, n_1457, n_1456);
not NOT1_3030 (n_1443, wire75);
and AND2_3031 (wire76, n_1405, n_1404);
or OR2_3032 (wire97, n_1405, n_1404);
not NOT1_3033 (n_1415, wire110);
and AND2_3034 (wire111, n_1366, n_1365);
or OR2_3035 (wire131, n_1366, n_1365);
and AND2_3036 (wire136, n_1342, n_1341);
not NOT1_3037 (n_1368, wire144);
not NOT1_3038 (n_1382, wire146);
or OR2_3039 (wire154, n_1342, n_1341);
or OR2_3040 (n_1352, wire166, n_1326);
not NOT1_3041 (n_1335, wire172);
not NOT1_3042 (n_1464, wire52);
or OR2_3043 (n_1483, wire62, n_1443);
or OR2_3044 (wire87, n_1415, n_1371);
or OR2_3045 (n_1430, wire88, n_1415);
not NOT1_3046 (n_1426, wire97);
or OR2_3047 (wire107, n_1368, n_1367);
and AND2_3048 (wire125, n_1352, n_1351);
and AND2_3049 (wire130, n_1368, n_1367);
not NOT1_3050 (n_1389, wire131);
or OR2_3051 (wire147, n_1352, n_1351);
not NOT1_3052 (n_1364, wire154);
or OR2_3053 (wire158, wire157, n_1335);
or OR2_3054 (n6170, wire42, n_1464);
or OR2_3055 (wire44, n_1464, n_1410);
and AND2_3056 (wire55, n_1431, n_1430);
or OR2_3057 (wire73, n_1431, n_1430);
or OR2_3058 (n_1438, wire76, n_1426);
or OR2_3059 (wire77, n_1426, n_1377);
not NOT1_3060 (n_1437, wire87);
or OR2_3061 (n_1407, wire111, n_1389);
not NOT1_3062 (n_1383, wire130);
or OR2_3063 (wire132, n_1364, n_1320);
or OR2_3064 (n_1381, wire136, n_1364);
not NOT1_3065 (n_1374, wire147);
not NOT1_3066 (n_1361, wire158);
not NOT1_3067 (n_1471, wire44);
and AND2_3068 (wire50, n_1438, n_1437);
or OR2_3069 (wire66, n_1438, n_1437);
and AND2_3070 (wire71, n_1407, n_1406);
not NOT1_3071 (n_1450, wire73);
not NOT1_3072 (n_1447, wire77);
or OR2_3073 (wire96, n_1407, n_1406);
and AND2_3074 (wire101, n_1382, n_1381);
and AND2_3075 (wire108, wire107, n_1383);
or OR2_3076 (wire114, n_1361, n_1360);
or OR2_3077 (wire119, n_1382, n_1381);
or OR2_3078 (wire123, n_1374, n_1326);
or OR2_3079 (n_1395, wire125, n_1374);
not NOT1_3080 (n_1396, wire132);
and AND2_3081 (wire139, n_1361, n_1360);
not NOT1_3082 (wire1678, n_1383);
and AND2_3083 (wire34, n_1471, n_1470);
or OR2_3084 (wire39, n_1471, n_1470);
or OR2_3085 (n_1487, wire55, n_1450);
not NOT1_3086 (n_1458, wire66);
and AND2_3087 (wire93, n_1396, n_1395);
not NOT1_3088 (n_1434, wire96);
or OR2_3089 (wire105, n_1396, n_1395);
not NOT1_3090 (n_1473, wire108);
not NOT1_3091 (n_1400, wire119);
not NOT1_3092 (n_1402, wire123);
not NOT1_3093 (n_1375, wire139);
or OR2_3094 (wire1679, wire1678, n_1354);
not NOT1_3095 (n_1477, wire39);
or OR2_3096 (n_1491, wire50, n_1458);
or OR2_3097 (wire70, n_1434, n_1389);
or OR2_3098 (n_1446, wire71, n_1434);
or OR2_3099 (n_1425, wire101, n_1400);
not NOT1_3100 (n_1411, wire105);
and AND2_3101 (wire115, wire114, n_1375);
not NOT1_3102 (n_1527, wire1679);
not NOT1_3103 (wire1680, n_1375);
or OR2_3104 (wire33, n_1477, n_1419);
or OR2_3105 (n6180, wire34, n_1477);
and AND2_3106 (wire46, n_1447, n_1446);
or OR2_3107 (wire58, n_1447, n_1446);
and AND2_3108 (wire60, n_1425, n_1424);
and AND2_3109 (wire63, n_1527, n528);
not NOT1_3110 (n_1452, wire70);
or OR2_3111 (wire78, n_1425, n_1424);
or OR2_3112 (wire82, wire81, n_1527);
or OR2_3113 (n_1433, wire93, n_1411);
not NOT1_3114 (n_1401, wire115);
or OR2_3115 (wire1681, wire1680, n_1335);
not NOT1_3116 (n_1480, wire33);
and AND2_3117 (wire56, n_1433, n_1432);
not NOT1_3118 (n_1461, wire58);
or OR2_3119 (wire72, n_1433, n_1432);
not NOT1_3120 (n_1444, wire78);
and AND2_3121 (wire79, n_1402, n_1401);
not NOT1_3122 (n_1442, wire82);
or OR2_3123 (wire100, n_1402, n_1401);
not NOT1_3124 (n_1528, wire1681);
and AND2_3125 (wire31, n_1480, n_1479);
or OR2_3126 (wire32, n_1480, n_1479);
or OR2_3127 (n_1495, wire46, n_1461);
or OR2_3128 (n_1451, wire60, n_1444);
or OR2_3129 (wire61, n_1444, n_1400);
or OR2_3130 (n_1519, wire63, n_1442);
and AND2_3131 (wire68, n_1417, n_1528);
not NOT1_3132 (n_1445, wire72);
or OR2_3133 (wire86, n_1417, n_1528);
not NOT1_3134 (n_1423, wire100);
not NOT1_3135 (n_1481, wire32);
and AND2_3136 (wire43, n_1452, n_1451);
or OR2_3137 (wire54, n_1452, n_1451);
or OR2_3138 (n_1459, wire56, n_1445);
or OR2_3139 (wire59, n_1445, n_1411);
not NOT1_3140 (n_1460, wire61);
or OR2_3141 (n_1440, wire79, n_1423);
not NOT1_3142 (n_1435, wire86);
or OR2_3143 (wire30, n_1481, n_1429);
or OR2_3144 (n6190, wire31, n_1481);
and AND2_3145 (wire40, n_1460, n_1459);
or OR2_3146 (wire49, n_1460, n_1459);
and AND2_3147 (wire51, n_1440, n_1439);
not NOT1_3148 (n_1465, wire54);
not NOT1_3149 (n_1463, wire59);
or OR2_3150 (wire65, n_1440, n_1439);
or OR2_3151 (wire69, wire68, n_1435);
not NOT1_3152 (n_1484, wire30);
or OR2_3153 (n_1499, wire43, n_1465);
not NOT1_3154 (n_1469, wire49);
not NOT1_3155 (n_1453, wire65);
not NOT1_3156 (n_1449, wire69);
and AND2_3157 (wire28, n_1484, n_1483);
or OR2_3158 (wire29, n_1484, n_1483);
or OR2_3159 (n_1503, wire40, n_1469);
or OR2_3160 (wire47, n_1449, n_1448);
or OR2_3161 (n_1462, wire51, n_1453);
or OR2_3162 (wire53, n_1453, n_1423);
and AND2_3163 (wire57, n_1449, n_1448);
not NOT1_3164 (n_1485, wire29);
and AND2_3165 (wire38, n_1463, n_1462);
or OR2_3166 (wire45, n_1463, n_1462);
not NOT1_3167 (n_1468, wire53);
not NOT1_3168 (n_1454, wire57);
or OR2_3169 (wire27, n_1485, n_1443);
or OR2_3170 (n6200, wire28, n_1485);
not NOT1_3171 (n_1472, wire45);
and AND2_3172 (wire48, wire47, n_1454);
not NOT1_3173 (wire1676, n_1454);
not NOT1_3174 (n_1488, wire27);
or OR2_3175 (n_1507, wire38, n_1472);
not NOT1_3176 (n_1467, wire48);
or OR2_3177 (wire1677, wire1676, n_1435);
and AND2_3178 (wire24, n_1488, n_1487);
or OR2_3179 (wire26, n_1488, n_1487);
and AND2_3180 (wire36, n_1468, n_1467);
or OR2_3181 (wire41, n_1468, n_1467);
not NOT1_3182 (n_1526, wire1677);
not NOT1_3183 (n_1489, wire26);
and AND2_3184 (wire35, n_1526, n_1473);
or OR2_3185 (wire37, n_1526, n_1473);
not NOT1_3186 (n_1475, wire41);
or OR2_3187 (n6210, wire24, n_1489);
or OR2_3188 (wire25, n_1489, n_1450);
or OR2_3189 (n_1511, wire36, n_1475);
not NOT1_3190 (n_1476, wire37);
not NOT1_3191 (n_1492, wire25);
or OR2_3192 (n_1515, wire35, n_1476);
and AND2_3193 (wire21, n_1492, n_1491);
or OR2_3194 (wire23, n_1492, n_1491);
not NOT1_3195 (n_1493, wire23);
or OR2_3196 (n6220, wire21, n_1493);
or OR2_3197 (wire22, n_1493, n_1458);
not NOT1_3198 (n_1496, wire22);
and AND2_3199 (wire18, n_1496, n_1495);
or OR2_3200 (wire20, n_1496, n_1495);
not NOT1_3201 (n_1497, wire20);
or OR2_3202 (n6230, wire18, n_1497);
or OR2_3203 (wire19, n_1497, n_1461);
not NOT1_3204 (n_1500, wire19);
and AND2_3205 (wire16, n_1500, n_1499);
or OR2_3206 (wire17, n_1500, n_1499);
not NOT1_3207 (n_1501, wire17);
or OR2_3208 (wire15, n_1501, n_1465);
or OR2_3209 (n6240, wire16, n_1501);
not NOT1_3210 (n_1504, wire15);
and AND2_3211 (wire12, n_1504, n_1503);
or OR2_3212 (wire14, n_1504, n_1503);
not NOT1_3213 (n_1505, wire14);
or OR2_3214 (n6250, wire12, n_1505);
or OR2_3215 (wire13, n_1505, n_1469);
not NOT1_3216 (n_1508, wire13);
and AND2_3217 (wire10, n_1508, n_1507);
or OR2_3218 (wire11, n_1508, n_1507);
not NOT1_3219 (n_1509, wire11);
or OR2_3220 (wire9, n_1509, n_1472);
or OR2_3221 (n6260, wire10, n_1509);
not NOT1_3222 (n_1512, wire9);
and AND2_3223 (wire6, n_1512, n_1511);
or OR2_3224 (wire8, n_1512, n_1511);
not NOT1_3225 (n_1513, wire8);
or OR2_3226 (n6270, wire6, n_1513);
or OR2_3227 (wire7, n_1513, n_1475);
not NOT1_3228 (n_1516, wire7);
and AND2_3229 (wire3, n_1516, n_1515);
or OR2_3230 (wire5, n_1516, n_1515);
not NOT1_3231 (n_1517, wire5);
or OR2_3232 (n6280, wire3, n_1517);
or OR2_3233 (wire4, n_1517, n_1476);
not NOT1_3234 (n_1520, wire4);
and AND2_3235 (wire1, n_1520, n_1519);
or OR2_3236 (wire2, n_1520, n_1519);
not NOT1_3237 (n_1521, wire2);
or OR2_3238 (wire0, n_1521, n_1442);
or OR2_3239 (n6288, wire1, n_1521);
not NOT1_3240 (n6287, wire0);

endmodule